
module INSTRMEM ( ADDR_RD, DATA_OUT );
  input [31:0] ADDR_RD;
  output [31:0] DATA_OUT;


endmodule


module DATAMEM ( RST, RE, WE, ADDR, DATA_IN, DATA_OUT );
  input [31:0] ADDR;
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT;
  input RST, RE, WE;


endmodule


module REG_BITS32_0 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1, n2, n3, n4;

  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n3), .Q(O[31]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n3), .Q(O[30]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n3), .Q(O[29]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n3), .Q(O[28]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n3), .Q(O[27]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n3), .Q(O[26]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n3), .Q(O[25]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n3), .Q(O[24]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n2), .Q(O[23]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n2), .Q(O[22]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n2), .Q(O[21]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n2), .Q(O[20]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n2), .Q(O[19]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n2), .Q(O[18]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n2), .Q(O[17]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n2), .Q(O[16]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n2), .Q(O[15]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n2), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n2), .Q(O[13]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n2), .Q(O[12]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  BUF_X1 U2 ( .A(n4), .Z(n1) );
  BUF_X1 U3 ( .A(n4), .Z(n2) );
  BUF_X1 U4 ( .A(n4), .Z(n3) );
  INV_X1 U5 ( .A(RST), .ZN(n4) );
endmodule


module ADDER_0_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238;

  AND2_X1 U2 ( .A1(n118), .A2(n100), .ZN(n117) );
  AND2_X1 U3 ( .A1(n160), .A2(n229), .ZN(SUM[0]) );
  AND4_X1 U4 ( .A1(n58), .A2(n53), .A3(n45), .A4(n47), .ZN(n2) );
  AND2_X1 U5 ( .A1(n104), .A2(n16), .ZN(n3) );
  AND2_X1 U6 ( .A1(n36), .A2(n39), .ZN(n4) );
  CLKBUF_X1 U7 ( .A(n103), .Z(n5) );
  AND4_X1 U8 ( .A1(n172), .A2(n173), .A3(n174), .A4(n175), .ZN(n6) );
  OAI21_X1 U9 ( .B1(n32), .B2(n85), .A(n86), .ZN(n7) );
  OAI21_X1 U10 ( .B1(n32), .B2(n85), .A(n86), .ZN(n8) );
  OAI21_X1 U11 ( .B1(n32), .B2(n85), .A(n86), .ZN(n77) );
  AND2_X2 U12 ( .A1(n103), .A2(n102), .ZN(n32) );
  AND2_X1 U13 ( .A1(n209), .A2(n210), .ZN(n9) );
  OAI21_X1 U14 ( .B1(n29), .B2(n129), .A(n131), .ZN(n10) );
  INV_X1 U15 ( .A(n23), .ZN(n11) );
  AND2_X1 U16 ( .A1(n227), .A2(n228), .ZN(n12) );
  NAND2_X1 U17 ( .A1(n105), .A2(n3), .ZN(n103) );
  OAI21_X1 U18 ( .B1(n117), .B2(n99), .A(n101), .ZN(n13) );
  AOI21_X1 U19 ( .B1(n133), .B2(n142), .A(n30), .ZN(n14) );
  OAI21_X1 U20 ( .B1(n9), .B2(n186), .A(n185), .ZN(n15) );
  AOI21_X1 U21 ( .B1(n17), .B2(n89), .A(n87), .ZN(n90) );
  NAND2_X1 U22 ( .A1(n16), .A2(n104), .ZN(n121) );
  AOI21_X1 U23 ( .B1(n16), .B2(n106), .A(n107), .ZN(n122) );
  INV_X1 U24 ( .A(n130), .ZN(n30) );
  OAI21_X1 U25 ( .B1(n167), .B2(n154), .A(n151), .ZN(n164) );
  OAI21_X1 U26 ( .B1(n224), .B2(n225), .A(n36), .ZN(n222) );
  AOI21_X1 U27 ( .B1(n87), .B2(n88), .A(n22), .ZN(n86) );
  AOI21_X1 U28 ( .B1(n155), .B2(n164), .A(n150), .ZN(n161) );
  OAI21_X1 U29 ( .B1(n117), .B2(n99), .A(n101), .ZN(n114) );
  NOR2_X1 U30 ( .A1(n146), .A2(n163), .ZN(n162) );
  NOR2_X1 U31 ( .A1(n92), .A2(n22), .ZN(n91) );
  NAND4_X1 U32 ( .A1(n156), .A2(n157), .A3(n155), .A4(n158), .ZN(n132) );
  AND4_X1 U33 ( .A1(n133), .A2(n134), .A3(n126), .A4(n135), .ZN(n16) );
  AND4_X1 U34 ( .A1(n108), .A2(n109), .A3(n96), .A4(n110), .ZN(n17) );
  NOR2_X1 U35 ( .A1(n94), .A2(n113), .ZN(n112) );
  NOR2_X1 U36 ( .A1(n124), .A2(n138), .ZN(n137) );
  NAND2_X1 U37 ( .A1(n56), .A2(n57), .ZN(n54) );
  NAND2_X1 U38 ( .A1(n226), .A2(n39), .ZN(n34) );
  NAND2_X1 U39 ( .A1(n170), .A2(n152), .ZN(n168) );
  NAND2_X1 U40 ( .A1(n23), .A2(n156), .ZN(n170) );
  NAND2_X1 U41 ( .A1(n165), .A2(n155), .ZN(n166) );
  NAND2_X1 U42 ( .A1(n217), .A2(n218), .ZN(n223) );
  AND2_X1 U43 ( .A1(n181), .A2(n179), .ZN(n203) );
  NAND2_X1 U44 ( .A1(n45), .A2(n44), .ZN(n49) );
  OAI21_X1 U45 ( .B1(n50), .B2(n51), .A(n52), .ZN(n46) );
  NAND2_X1 U46 ( .A1(n65), .A2(n64), .ZN(n79) );
  NAND2_X1 U47 ( .A1(n73), .A2(n71), .ZN(n74) );
  NAND2_X1 U48 ( .A1(n43), .A2(n44), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n45), .A2(n46), .ZN(n43) );
  NAND2_X1 U50 ( .A1(n221), .A2(n217), .ZN(n220) );
  NAND2_X1 U51 ( .A1(n218), .A2(n222), .ZN(n221) );
  NAND2_X1 U52 ( .A1(n130), .A2(n133), .ZN(n143) );
  NAND2_X1 U53 ( .A1(n47), .A2(n48), .ZN(n41) );
  NAND2_X1 U54 ( .A1(n53), .A2(n52), .ZN(n55) );
  NAND2_X1 U55 ( .A1(n35), .A2(n36), .ZN(n33) );
  AND2_X1 U56 ( .A1(n101), .A2(n109), .ZN(n18) );
  AND2_X1 U57 ( .A1(n131), .A2(n134), .ZN(n19) );
  NAND2_X1 U58 ( .A1(n195), .A2(n216), .ZN(n219) );
  NAND2_X1 U59 ( .A1(n157), .A2(n151), .ZN(n169) );
  NAND2_X1 U60 ( .A1(n82), .A2(n81), .ZN(n159) );
  NAND2_X1 U61 ( .A1(n115), .A2(n96), .ZN(n116) );
  NAND2_X1 U62 ( .A1(n140), .A2(n126), .ZN(n141) );
  NAND2_X1 U63 ( .A1(n57), .A2(n58), .ZN(n59) );
  NAND2_X1 U64 ( .A1(n100), .A2(n108), .ZN(n120) );
  NAND2_X1 U65 ( .A1(n76), .A2(n78), .ZN(n84) );
  NAND2_X1 U66 ( .A1(n39), .A2(n40), .ZN(n37) );
  NAND2_X1 U67 ( .A1(n210), .A2(n200), .ZN(n212) );
  NAND2_X1 U68 ( .A1(n156), .A2(n152), .ZN(n171) );
  NAND2_X1 U69 ( .A1(n67), .A2(n68), .ZN(n60) );
  NAND2_X1 U70 ( .A1(n201), .A2(n185), .ZN(n208) );
  AND2_X1 U71 ( .A1(n67), .A2(n192), .ZN(n20) );
  AND2_X1 U72 ( .A1(n68), .A2(n64), .ZN(n232) );
  OAI21_X1 U73 ( .B1(n145), .B2(n146), .A(n147), .ZN(n106) );
  AOI21_X1 U74 ( .B1(n148), .B2(n149), .A(n150), .ZN(n145) );
  NAND2_X1 U75 ( .A1(n151), .A2(n152), .ZN(n149) );
  OAI21_X1 U76 ( .B1(n93), .B2(n94), .A(n95), .ZN(n87) );
  AOI21_X1 U77 ( .B1(n96), .B2(n97), .A(n98), .ZN(n93) );
  OAI21_X1 U78 ( .B1(n99), .B2(n100), .A(n101), .ZN(n97) );
  OAI21_X1 U79 ( .B1(n123), .B2(n124), .A(n125), .ZN(n107) );
  AOI21_X1 U80 ( .B1(n126), .B2(n127), .A(n128), .ZN(n123) );
  OAI21_X1 U81 ( .B1(n129), .B2(n130), .A(n131), .ZN(n127) );
  OAI21_X1 U82 ( .B1(n4), .B2(n214), .A(n215), .ZN(n197) );
  AND2_X1 U83 ( .A1(n216), .A2(n217), .ZN(n215) );
  NAND2_X1 U84 ( .A1(n218), .A2(n35), .ZN(n214) );
  AND2_X1 U85 ( .A1(n48), .A2(n44), .ZN(n235) );
  NAND2_X1 U86 ( .A1(n238), .A2(n45), .ZN(n234) );
  NAND2_X1 U87 ( .A1(n80), .A2(n81), .ZN(n66) );
  NAND2_X1 U88 ( .A1(n82), .A2(n83), .ZN(n80) );
  INV_X1 U89 ( .A(n160), .ZN(n83) );
  NAND2_X1 U90 ( .A1(n184), .A2(n185), .ZN(n183) );
  INV_X1 U91 ( .A(n176), .ZN(n175) );
  OAI21_X1 U92 ( .B1(n177), .B2(n178), .A(n179), .ZN(n176) );
  NOR2_X1 U93 ( .A1(n182), .A2(n183), .ZN(n177) );
  OR2_X1 U94 ( .A1(B[20]), .A2(A[20]), .ZN(n133) );
  OR2_X1 U95 ( .A1(B[6]), .A2(A[6]), .ZN(n45) );
  OR2_X1 U96 ( .A1(B[14]), .A2(A[14]), .ZN(n180) );
  OR2_X1 U97 ( .A1(B[18]), .A2(A[18]), .ZN(n155) );
  OR2_X1 U98 ( .A1(B[22]), .A2(A[22]), .ZN(n126) );
  OR2_X1 U99 ( .A1(B[26]), .A2(A[26]), .ZN(n96) );
  NAND2_X1 U100 ( .A1(B[0]), .A2(A[0]), .ZN(n231) );
  OR2_X1 U101 ( .A1(B[7]), .A2(A[7]), .ZN(n47) );
  OR2_X1 U102 ( .A1(B[5]), .A2(A[5]), .ZN(n53) );
  OR2_X1 U103 ( .A1(B[9]), .A2(A[9]), .ZN(n35) );
  OR2_X1 U104 ( .A1(B[16]), .A2(A[16]), .ZN(n156) );
  OR2_X1 U105 ( .A1(B[4]), .A2(A[4]), .ZN(n58) );
  OR2_X1 U106 ( .A1(B[21]), .A2(A[21]), .ZN(n134) );
  OR2_X1 U107 ( .A1(B[25]), .A2(A[25]), .ZN(n109) );
  OR2_X1 U108 ( .A1(B[11]), .A2(A[11]), .ZN(n195) );
  OR2_X1 U109 ( .A1(B[24]), .A2(A[24]), .ZN(n108) );
  OR2_X1 U110 ( .A1(B[1]), .A2(A[1]), .ZN(n82) );
  NAND2_X1 U111 ( .A1(B[2]), .A2(A[2]), .ZN(n64) );
  OR2_X1 U112 ( .A1(B[28]), .A2(A[28]), .ZN(n88) );
  OR2_X1 U113 ( .A1(B[29]), .A2(A[29]), .ZN(n78) );
  OR2_X1 U114 ( .A1(B[8]), .A2(A[8]), .ZN(n40) );
  OR2_X1 U115 ( .A1(B[12]), .A2(A[12]), .ZN(n200) );
  OR2_X1 U116 ( .A1(B[3]), .A2(A[3]), .ZN(n67) );
  OR2_X1 U117 ( .A1(B[13]), .A2(A[13]), .ZN(n201) );
  OR2_X1 U118 ( .A1(B[19]), .A2(A[19]), .ZN(n158) );
  OR2_X1 U119 ( .A1(B[23]), .A2(A[23]), .ZN(n135) );
  OR2_X1 U120 ( .A1(B[27]), .A2(A[27]), .ZN(n110) );
  OR2_X1 U121 ( .A1(B[15]), .A2(A[15]), .ZN(n181) );
  OR2_X1 U122 ( .A1(B[30]), .A2(A[30]), .ZN(n71) );
  OR2_X1 U123 ( .A1(B[0]), .A2(A[0]), .ZN(n229) );
  OR2_X1 U124 ( .A1(B[10]), .A2(A[10]), .ZN(n218) );
  OR2_X1 U125 ( .A1(B[17]), .A2(A[17]), .ZN(n157) );
  XOR2_X1 U126 ( .A(B[31]), .B(A[31]), .Z(n21) );
  NAND2_X1 U127 ( .A1(B[20]), .A2(A[20]), .ZN(n130) );
  AND2_X1 U128 ( .A1(B[28]), .A2(A[28]), .ZN(n22) );
  NAND2_X1 U129 ( .A1(B[16]), .A2(A[16]), .ZN(n152) );
  NAND2_X1 U130 ( .A1(B[8]), .A2(A[8]), .ZN(n39) );
  NAND2_X1 U131 ( .A1(B[9]), .A2(A[9]), .ZN(n36) );
  NAND2_X1 U132 ( .A1(B[17]), .A2(A[17]), .ZN(n151) );
  NAND2_X1 U133 ( .A1(B[25]), .A2(A[25]), .ZN(n101) );
  NAND2_X1 U134 ( .A1(B[6]), .A2(A[6]), .ZN(n44) );
  NAND2_X1 U135 ( .A1(B[13]), .A2(A[13]), .ZN(n185) );
  OR2_X1 U136 ( .A1(B[2]), .A2(A[2]), .ZN(n65) );
  NAND2_X1 U137 ( .A1(B[5]), .A2(A[5]), .ZN(n52) );
  NAND2_X1 U138 ( .A1(B[10]), .A2(A[10]), .ZN(n217) );
  NAND2_X1 U139 ( .A1(B[4]), .A2(A[4]), .ZN(n57) );
  NAND2_X1 U140 ( .A1(B[21]), .A2(A[21]), .ZN(n131) );
  NAND2_X1 U141 ( .A1(B[24]), .A2(A[24]), .ZN(n100) );
  NAND2_X1 U142 ( .A1(B[1]), .A2(A[1]), .ZN(n81) );
  NAND2_X1 U143 ( .A1(B[14]), .A2(A[14]), .ZN(n184) );
  NAND2_X1 U144 ( .A1(B[29]), .A2(A[29]), .ZN(n76) );
  NAND2_X1 U145 ( .A1(B[0]), .A2(A[0]), .ZN(n160) );
  NAND2_X1 U146 ( .A1(B[3]), .A2(A[3]), .ZN(n68) );
  NAND2_X1 U147 ( .A1(B[7]), .A2(A[7]), .ZN(n48) );
  NAND2_X1 U148 ( .A1(B[11]), .A2(A[11]), .ZN(n216) );
  NAND2_X1 U149 ( .A1(B[23]), .A2(A[23]), .ZN(n125) );
  NAND2_X1 U150 ( .A1(B[15]), .A2(A[15]), .ZN(n179) );
  NAND2_X1 U151 ( .A1(B[19]), .A2(A[19]), .ZN(n147) );
  NAND2_X1 U152 ( .A1(B[27]), .A2(A[27]), .ZN(n95) );
  NAND2_X1 U153 ( .A1(B[22]), .A2(A[22]), .ZN(n140) );
  NAND2_X1 U154 ( .A1(B[18]), .A2(A[18]), .ZN(n165) );
  NAND2_X1 U155 ( .A1(B[26]), .A2(A[26]), .ZN(n115) );
  NAND2_X1 U156 ( .A1(B[30]), .A2(A[30]), .ZN(n73) );
  NAND2_X1 U157 ( .A1(B[12]), .A2(A[12]), .ZN(n210) );
  XNOR2_X1 U158 ( .A(n49), .B(n46), .ZN(SUM[6]) );
  XNOR2_X1 U159 ( .A(n223), .B(n222), .ZN(SUM[10]) );
  XNOR2_X1 U160 ( .A(n166), .B(n164), .ZN(SUM[18]) );
  XNOR2_X1 U161 ( .A(n74), .B(n31), .ZN(SUM[30]) );
  XNOR2_X1 U162 ( .A(n33), .B(n34), .ZN(SUM[9]) );
  XNOR2_X1 U163 ( .A(n55), .B(n54), .ZN(SUM[5]) );
  XNOR2_X1 U164 ( .A(n169), .B(n168), .ZN(SUM[17]) );
  XNOR2_X1 U165 ( .A(n219), .B(n220), .ZN(SUM[11]) );
  XNOR2_X1 U166 ( .A(n41), .B(n42), .ZN(SUM[7]) );
  XNOR2_X1 U167 ( .A(n161), .B(n162), .ZN(SUM[19]) );
  XNOR2_X1 U168 ( .A(n90), .B(n91), .ZN(SUM[28]) );
  XNOR2_X1 U169 ( .A(n79), .B(n66), .ZN(SUM[2]) );
  XNOR2_X1 U170 ( .A(n159), .B(n83), .ZN(SUM[1]) );
  XNOR2_X1 U171 ( .A(n208), .B(n207), .ZN(SUM[13]) );
  NAND2_X1 U172 ( .A1(n180), .A2(n181), .ZN(n178) );
  NAND2_X1 U173 ( .A1(n180), .A2(n184), .ZN(n206) );
  NOR2_X1 U174 ( .A1(n188), .A2(n194), .ZN(n191) );
  NAND2_X1 U175 ( .A1(n209), .A2(n210), .ZN(n207) );
  NAND4_X1 U176 ( .A1(n200), .A2(n201), .A3(n180), .A4(n181), .ZN(n189) );
  OAI21_X1 U177 ( .B1(n12), .B2(n24), .A(n213), .ZN(n211) );
  OAI21_X1 U178 ( .B1(n9), .B2(n186), .A(n185), .ZN(n204) );
  NAND4_X1 U179 ( .A1(n58), .A2(n53), .A3(n45), .A4(n47), .ZN(n188) );
  NAND4_X1 U180 ( .A1(n173), .A2(n174), .A3(n172), .A4(n175), .ZN(n23) );
  NAND4_X1 U181 ( .A1(n172), .A2(n173), .A3(n174), .A4(n175), .ZN(n105) );
  INV_X1 U182 ( .A(n198), .ZN(n24) );
  NAND4_X1 U183 ( .A1(n195), .A2(n218), .A3(n35), .A4(n40), .ZN(n190) );
  OAI21_X1 U184 ( .B1(n14), .B2(n129), .A(n131), .ZN(n139) );
  CLKBUF_X1 U185 ( .A(n117), .Z(n25) );
  CLKBUF_X1 U186 ( .A(n20), .Z(n26) );
  XNOR2_X1 U187 ( .A(n84), .B(n8), .ZN(SUM[29]) );
  AOI21_X1 U188 ( .B1(n70), .B2(n71), .A(n72), .ZN(n69) );
  NAND2_X1 U189 ( .A1(n7), .A2(n78), .ZN(n27) );
  OAI21_X1 U190 ( .B1(n11), .B2(n121), .A(n122), .ZN(n28) );
  NAND2_X1 U191 ( .A1(n38), .A2(n40), .ZN(n226) );
  XNOR2_X1 U192 ( .A(n37), .B(n38), .ZN(SUM[8]) );
  NAND2_X1 U193 ( .A1(n227), .A2(n228), .ZN(n38) );
  NAND2_X1 U194 ( .A1(n82), .A2(n65), .ZN(n230) );
  AOI21_X1 U195 ( .B1(n133), .B2(n142), .A(n30), .ZN(n29) );
  XNOR2_X1 U196 ( .A(n111), .B(n112), .ZN(SUM[27]) );
  NAND2_X1 U197 ( .A1(n27), .A2(n76), .ZN(n31) );
  NAND2_X1 U198 ( .A1(n75), .A2(n76), .ZN(n70) );
  NAND2_X1 U199 ( .A1(n77), .A2(n78), .ZN(n75) );
  OAI21_X1 U200 ( .B1(n6), .B2(n132), .A(n144), .ZN(n142) );
  OAI21_X1 U201 ( .B1(n6), .B2(n121), .A(n122), .ZN(n119) );
  NAND2_X1 U202 ( .A1(n119), .A2(n108), .ZN(n118) );
  AOI21_X1 U203 ( .B1(n13), .B2(n96), .A(n98), .ZN(n111) );
  OAI211_X1 U204 ( .C1(n230), .C2(n231), .A(n232), .B(n233), .ZN(n192) );
  XNOR2_X1 U205 ( .A(n202), .B(n203), .ZN(SUM[15]) );
  AOI21_X1 U206 ( .B1(n16), .B2(n106), .A(n107), .ZN(n102) );
  NOR2_X1 U207 ( .A1(n189), .A2(n190), .ZN(n193) );
  NAND2_X1 U208 ( .A1(n102), .A2(n5), .ZN(n89) );
  XNOR2_X1 U209 ( .A(n206), .B(n204), .ZN(SUM[14]) );
  XNOR2_X1 U210 ( .A(n212), .B(n211), .ZN(SUM[12]) );
  XNOR2_X1 U211 ( .A(n59), .B(n26), .ZN(SUM[4]) );
  AOI21_X1 U212 ( .B1(n15), .B2(n180), .A(n205), .ZN(n202) );
  NAND2_X1 U213 ( .A1(n211), .A2(n200), .ZN(n209) );
  NAND2_X1 U214 ( .A1(n26), .A2(n58), .ZN(n56) );
  NAND2_X1 U215 ( .A1(n2), .A2(n20), .ZN(n228) );
  XNOR2_X1 U216 ( .A(n69), .B(n21), .ZN(SUM[31]) );
  XNOR2_X1 U217 ( .A(n136), .B(n137), .ZN(SUM[23]) );
  AOI21_X1 U218 ( .B1(n139), .B2(n126), .A(n128), .ZN(n136) );
  INV_X1 U219 ( .A(n53), .ZN(n51) );
  INV_X1 U220 ( .A(n54), .ZN(n50) );
  XNOR2_X1 U221 ( .A(n60), .B(n61), .ZN(SUM[3]) );
  OAI21_X1 U222 ( .B1(n62), .B2(n63), .A(n64), .ZN(n61) );
  INV_X1 U223 ( .A(n65), .ZN(n63) );
  INV_X1 U224 ( .A(n66), .ZN(n62) );
  INV_X1 U225 ( .A(n73), .ZN(n72) );
  NAND2_X1 U226 ( .A1(n17), .A2(n88), .ZN(n85) );
  INV_X1 U227 ( .A(n88), .ZN(n92) );
  INV_X1 U228 ( .A(n95), .ZN(n113) );
  INV_X1 U229 ( .A(n110), .ZN(n94) );
  INV_X1 U230 ( .A(n115), .ZN(n98) );
  XNOR2_X1 U231 ( .A(n116), .B(n114), .ZN(SUM[26]) );
  INV_X1 U232 ( .A(n109), .ZN(n99) );
  XNOR2_X1 U233 ( .A(n25), .B(n18), .ZN(SUM[25]) );
  XNOR2_X1 U234 ( .A(n120), .B(n28), .ZN(SUM[24]) );
  INV_X1 U235 ( .A(n132), .ZN(n104) );
  INV_X1 U236 ( .A(n125), .ZN(n138) );
  INV_X1 U237 ( .A(n135), .ZN(n124) );
  INV_X1 U238 ( .A(n140), .ZN(n128) );
  XNOR2_X1 U239 ( .A(n10), .B(n141), .ZN(SUM[22]) );
  INV_X1 U240 ( .A(n134), .ZN(n129) );
  XNOR2_X1 U241 ( .A(n29), .B(n19), .ZN(SUM[21]) );
  XNOR2_X1 U242 ( .A(n143), .B(n142), .ZN(SUM[20]) );
  INV_X1 U243 ( .A(n106), .ZN(n144) );
  NOR2_X1 U244 ( .A1(n153), .A2(n154), .ZN(n148) );
  INV_X1 U245 ( .A(n155), .ZN(n153) );
  INV_X1 U246 ( .A(n147), .ZN(n163) );
  INV_X1 U247 ( .A(n158), .ZN(n146) );
  INV_X1 U248 ( .A(n165), .ZN(n150) );
  INV_X1 U249 ( .A(n157), .ZN(n154) );
  INV_X1 U250 ( .A(n168), .ZN(n167) );
  XNOR2_X1 U251 ( .A(n171), .B(n23), .ZN(SUM[16]) );
  NOR2_X1 U252 ( .A1(n186), .A2(n187), .ZN(n182) );
  NAND2_X1 U253 ( .A1(A[12]), .A2(B[12]), .ZN(n187) );
  NAND3_X1 U254 ( .A1(n191), .A2(n193), .A3(n192), .ZN(n174) );
  NAND3_X1 U255 ( .A1(n195), .A2(n196), .A3(n197), .ZN(n173) );
  NAND4_X1 U256 ( .A1(n198), .A2(n196), .A3(n47), .A4(n199), .ZN(n172) );
  INV_X1 U257 ( .A(n189), .ZN(n196) );
  INV_X1 U258 ( .A(n190), .ZN(n198) );
  INV_X1 U259 ( .A(n184), .ZN(n205) );
  INV_X1 U260 ( .A(n201), .ZN(n186) );
  NAND2_X1 U261 ( .A1(n195), .A2(n197), .ZN(n213) );
  INV_X1 U262 ( .A(n35), .ZN(n225) );
  INV_X1 U263 ( .A(n34), .ZN(n224) );
  INV_X1 U264 ( .A(n67), .ZN(n194) );
  NAND3_X1 U265 ( .A1(A[1]), .A2(B[1]), .A3(n65), .ZN(n233) );
  NAND2_X1 U266 ( .A1(n47), .A2(n199), .ZN(n227) );
  NAND3_X1 U267 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n199) );
  NAND3_X1 U268 ( .A1(n53), .A2(n45), .A3(n237), .ZN(n236) );
  INV_X1 U269 ( .A(n57), .ZN(n237) );
  INV_X1 U270 ( .A(n52), .ZN(n238) );
endmodule


module ADDER_0 ( A, B, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;


  ADDER_0_DW01_add_2 add_16 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module MUX21_NBIT5_0 ( IN0, IN1, S, O );
  input [4:0] IN0;
  input [4:0] IN1;
  output [4:0] O;
  input S;
  wire   n7, n8, n9, n10, n11, n6;

  INV_X1 U1 ( .A(n8), .ZN(O[3]) );
  AOI22_X1 U2 ( .A1(IN0[3]), .A2(n6), .B1(IN1[3]), .B2(S), .ZN(n8) );
  INV_X1 U3 ( .A(n11), .ZN(O[0]) );
  AOI22_X1 U4 ( .A1(IN0[0]), .A2(n6), .B1(IN1[0]), .B2(S), .ZN(n11) );
  INV_X1 U5 ( .A(n9), .ZN(O[2]) );
  AOI22_X1 U6 ( .A1(IN0[2]), .A2(n6), .B1(IN1[2]), .B2(S), .ZN(n9) );
  INV_X1 U7 ( .A(n10), .ZN(O[1]) );
  AOI22_X1 U8 ( .A1(IN0[1]), .A2(n6), .B1(IN1[1]), .B2(S), .ZN(n10) );
  INV_X1 U9 ( .A(n7), .ZN(O[4]) );
  AOI22_X1 U10 ( .A1(IN0[4]), .A2(n6), .B1(S), .B2(IN1[4]), .ZN(n7) );
  INV_X1 U11 ( .A(S), .ZN(n6) );
endmodule


module MUX21_NBIT32_0 ( IN0, IN1, S, O );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] O;
  input S;
  wire   n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n1, n2, n3, n68;

  BUF_X1 U1 ( .A(n68), .Z(n1) );
  BUF_X1 U2 ( .A(n68), .Z(n2) );
  BUF_X1 U3 ( .A(n68), .Z(n3) );
  INV_X1 U4 ( .A(n53), .ZN(O[20]) );
  AOI22_X1 U5 ( .A1(IN0[20]), .A2(n2), .B1(IN1[20]), .B2(S), .ZN(n53) );
  INV_X1 U6 ( .A(n52), .ZN(O[21]) );
  AOI22_X1 U7 ( .A1(IN0[21]), .A2(n2), .B1(IN1[21]), .B2(S), .ZN(n52) );
  INV_X1 U8 ( .A(n51), .ZN(O[22]) );
  AOI22_X1 U9 ( .A1(IN0[22]), .A2(n2), .B1(IN1[22]), .B2(S), .ZN(n51) );
  INV_X1 U10 ( .A(n50), .ZN(O[23]) );
  AOI22_X1 U11 ( .A1(IN0[23]), .A2(n2), .B1(IN1[23]), .B2(S), .ZN(n50) );
  INV_X1 U12 ( .A(n49), .ZN(O[24]) );
  AOI22_X1 U13 ( .A1(IN0[24]), .A2(n2), .B1(IN1[24]), .B2(S), .ZN(n49) );
  INV_X1 U14 ( .A(n48), .ZN(O[25]) );
  AOI22_X1 U15 ( .A1(IN0[25]), .A2(n2), .B1(IN1[25]), .B2(S), .ZN(n48) );
  INV_X1 U16 ( .A(n47), .ZN(O[26]) );
  AOI22_X1 U17 ( .A1(IN0[26]), .A2(n2), .B1(IN1[26]), .B2(S), .ZN(n47) );
  INV_X1 U18 ( .A(n46), .ZN(O[27]) );
  AOI22_X1 U19 ( .A1(IN0[27]), .A2(n2), .B1(IN1[27]), .B2(S), .ZN(n46) );
  INV_X1 U20 ( .A(n45), .ZN(O[28]) );
  AOI22_X1 U21 ( .A1(IN0[28]), .A2(n2), .B1(IN1[28]), .B2(S), .ZN(n45) );
  INV_X1 U22 ( .A(n44), .ZN(O[29]) );
  AOI22_X1 U23 ( .A1(IN0[29]), .A2(n2), .B1(IN1[29]), .B2(S), .ZN(n44) );
  INV_X1 U24 ( .A(n42), .ZN(O[30]) );
  AOI22_X1 U25 ( .A1(IN0[30]), .A2(n2), .B1(IN1[30]), .B2(S), .ZN(n42) );
  INV_X1 U26 ( .A(n41), .ZN(O[31]) );
  AOI22_X1 U27 ( .A1(IN0[31]), .A2(n3), .B1(IN1[31]), .B2(S), .ZN(n41) );
  INV_X1 U28 ( .A(n35), .ZN(O[8]) );
  AOI22_X1 U29 ( .A1(IN0[8]), .A2(n3), .B1(IN1[8]), .B2(S), .ZN(n35) );
  INV_X1 U30 ( .A(n34), .ZN(O[9]) );
  AOI22_X1 U31 ( .A1(IN0[9]), .A2(n3), .B1(S), .B2(IN1[9]), .ZN(n34) );
  INV_X1 U32 ( .A(n64), .ZN(O[10]) );
  AOI22_X1 U33 ( .A1(IN0[10]), .A2(n1), .B1(IN1[10]), .B2(S), .ZN(n64) );
  INV_X1 U34 ( .A(n63), .ZN(O[11]) );
  AOI22_X1 U35 ( .A1(IN0[11]), .A2(n1), .B1(IN1[11]), .B2(S), .ZN(n63) );
  INV_X1 U36 ( .A(n62), .ZN(O[12]) );
  AOI22_X1 U37 ( .A1(IN0[12]), .A2(n1), .B1(IN1[12]), .B2(S), .ZN(n62) );
  INV_X1 U38 ( .A(n61), .ZN(O[13]) );
  AOI22_X1 U39 ( .A1(IN0[13]), .A2(n1), .B1(IN1[13]), .B2(S), .ZN(n61) );
  INV_X1 U40 ( .A(n60), .ZN(O[14]) );
  AOI22_X1 U41 ( .A1(IN0[14]), .A2(n1), .B1(IN1[14]), .B2(S), .ZN(n60) );
  INV_X1 U42 ( .A(n59), .ZN(O[15]) );
  AOI22_X1 U43 ( .A1(IN0[15]), .A2(n1), .B1(IN1[15]), .B2(S), .ZN(n59) );
  INV_X1 U44 ( .A(n58), .ZN(O[16]) );
  AOI22_X1 U45 ( .A1(IN0[16]), .A2(n1), .B1(IN1[16]), .B2(S), .ZN(n58) );
  INV_X1 U46 ( .A(n57), .ZN(O[17]) );
  AOI22_X1 U47 ( .A1(IN0[17]), .A2(n1), .B1(IN1[17]), .B2(S), .ZN(n57) );
  INV_X1 U48 ( .A(n56), .ZN(O[18]) );
  AOI22_X1 U49 ( .A1(IN0[18]), .A2(n1), .B1(IN1[18]), .B2(S), .ZN(n56) );
  INV_X1 U50 ( .A(n55), .ZN(O[19]) );
  AOI22_X1 U51 ( .A1(IN0[19]), .A2(n1), .B1(IN1[19]), .B2(S), .ZN(n55) );
  INV_X1 U52 ( .A(n65), .ZN(O[0]) );
  AOI22_X1 U53 ( .A1(IN0[0]), .A2(n1), .B1(IN1[0]), .B2(S), .ZN(n65) );
  INV_X1 U54 ( .A(n54), .ZN(O[1]) );
  AOI22_X1 U55 ( .A1(IN0[1]), .A2(n1), .B1(IN1[1]), .B2(S), .ZN(n54) );
  INV_X1 U56 ( .A(n43), .ZN(O[2]) );
  AOI22_X1 U57 ( .A1(IN0[2]), .A2(n2), .B1(IN1[2]), .B2(S), .ZN(n43) );
  INV_X1 U58 ( .A(n40), .ZN(O[3]) );
  AOI22_X1 U59 ( .A1(IN0[3]), .A2(n3), .B1(IN1[3]), .B2(S), .ZN(n40) );
  INV_X1 U60 ( .A(n39), .ZN(O[4]) );
  AOI22_X1 U61 ( .A1(IN0[4]), .A2(n3), .B1(IN1[4]), .B2(S), .ZN(n39) );
  INV_X1 U62 ( .A(n38), .ZN(O[5]) );
  AOI22_X1 U63 ( .A1(IN0[5]), .A2(n3), .B1(IN1[5]), .B2(S), .ZN(n38) );
  INV_X1 U64 ( .A(n37), .ZN(O[6]) );
  AOI22_X1 U65 ( .A1(IN0[6]), .A2(n3), .B1(IN1[6]), .B2(S), .ZN(n37) );
  INV_X1 U66 ( .A(n36), .ZN(O[7]) );
  AOI22_X1 U67 ( .A1(IN0[7]), .A2(n3), .B1(IN1[7]), .B2(S), .ZN(n36) );
  INV_X1 U68 ( .A(S), .ZN(n68) );
endmodule


module MUX21_NBIT5_1 ( IN0, IN1, S, O );
  input [4:0] IN0;
  input [4:0] IN1;
  output [4:0] O;
  input S;
  wire   n6, n12, n13, n14, n15, n16;

  INV_X1 U1 ( .A(n14), .ZN(O[2]) );
  AOI22_X1 U2 ( .A1(IN0[2]), .A2(n6), .B1(IN1[2]), .B2(S), .ZN(n14) );
  INV_X1 U3 ( .A(n13), .ZN(O[1]) );
  AOI22_X1 U4 ( .A1(IN0[1]), .A2(n6), .B1(IN1[1]), .B2(S), .ZN(n13) );
  INV_X1 U5 ( .A(n12), .ZN(O[0]) );
  AOI22_X1 U6 ( .A1(IN0[0]), .A2(n6), .B1(IN1[0]), .B2(S), .ZN(n12) );
  INV_X1 U7 ( .A(n16), .ZN(O[4]) );
  AOI22_X1 U8 ( .A1(IN0[4]), .A2(n6), .B1(S), .B2(IN1[4]), .ZN(n16) );
  INV_X1 U9 ( .A(n15), .ZN(O[3]) );
  AOI22_X1 U10 ( .A1(IN0[3]), .A2(n6), .B1(IN1[3]), .B2(S), .ZN(n15) );
  INV_X1 U11 ( .A(S), .ZN(n6) );
endmodule


module RF ( RST, WE, ADDR_RD1, ADDR_RD2, ADDR_WR, DATA_IN, DATA_OUT1, 
        DATA_OUT2 );
  input [4:0] ADDR_RD1;
  input [4:0] ADDR_RD2;
  input [4:0] ADDR_WR;
  input [31:0] DATA_IN;
  output [31:0] DATA_OUT1;
  output [31:0] DATA_OUT2;
  input RST, WE;
  wire   \REGS[0][31] , \REGS[0][30] , \REGS[0][29] , \REGS[0][28] ,
         \REGS[0][27] , \REGS[0][26] , \REGS[0][25] , \REGS[0][24] ,
         \REGS[0][23] , \REGS[0][22] , \REGS[0][21] , \REGS[0][20] ,
         \REGS[0][19] , \REGS[0][18] , \REGS[0][17] , \REGS[0][16] ,
         \REGS[0][15] , \REGS[0][14] , \REGS[0][13] , \REGS[0][12] ,
         \REGS[0][11] , \REGS[0][10] , \REGS[0][9] , \REGS[0][8] ,
         \REGS[0][7] , \REGS[0][6] , \REGS[0][5] , \REGS[0][4] , \REGS[0][3] ,
         \REGS[0][2] , \REGS[0][1] , \REGS[0][0] , \REGS[1][31] ,
         \REGS[1][30] , \REGS[1][29] , \REGS[1][28] , \REGS[1][27] ,
         \REGS[1][26] , \REGS[1][25] , \REGS[1][24] , \REGS[1][23] ,
         \REGS[1][22] , \REGS[1][21] , \REGS[1][20] , \REGS[1][19] ,
         \REGS[1][18] , \REGS[1][17] , \REGS[1][16] , \REGS[1][15] ,
         \REGS[1][14] , \REGS[1][13] , \REGS[1][12] , \REGS[1][11] ,
         \REGS[1][10] , \REGS[1][9] , \REGS[1][8] , \REGS[1][7] , \REGS[1][6] ,
         \REGS[1][5] , \REGS[1][4] , \REGS[1][3] , \REGS[1][2] , \REGS[1][1] ,
         \REGS[1][0] , \REGS[2][31] , \REGS[2][30] , \REGS[2][29] ,
         \REGS[2][28] , \REGS[2][27] , \REGS[2][26] , \REGS[2][25] ,
         \REGS[2][24] , \REGS[2][23] , \REGS[2][22] , \REGS[2][21] ,
         \REGS[2][20] , \REGS[2][19] , \REGS[2][18] , \REGS[2][17] ,
         \REGS[2][16] , \REGS[2][15] , \REGS[2][14] , \REGS[2][13] ,
         \REGS[2][12] , \REGS[2][11] , \REGS[2][10] , \REGS[2][9] ,
         \REGS[2][8] , \REGS[2][7] , \REGS[2][6] , \REGS[2][5] , \REGS[2][4] ,
         \REGS[2][3] , \REGS[2][2] , \REGS[2][1] , \REGS[2][0] , \REGS[3][31] ,
         \REGS[3][30] , \REGS[3][29] , \REGS[3][28] , \REGS[3][27] ,
         \REGS[3][26] , \REGS[3][25] , \REGS[3][24] , \REGS[3][23] ,
         \REGS[3][22] , \REGS[3][21] , \REGS[3][20] , \REGS[3][19] ,
         \REGS[3][18] , \REGS[3][17] , \REGS[3][16] , \REGS[3][15] ,
         \REGS[3][14] , \REGS[3][13] , \REGS[3][12] , \REGS[3][11] ,
         \REGS[3][10] , \REGS[3][9] , \REGS[3][8] , \REGS[3][7] , \REGS[3][6] ,
         \REGS[3][5] , \REGS[3][4] , \REGS[3][3] , \REGS[3][2] , \REGS[3][1] ,
         \REGS[3][0] , \REGS[4][31] , \REGS[4][30] , \REGS[4][29] ,
         \REGS[4][28] , \REGS[4][27] , \REGS[4][26] , \REGS[4][25] ,
         \REGS[4][24] , \REGS[4][23] , \REGS[4][22] , \REGS[4][21] ,
         \REGS[4][20] , \REGS[4][19] , \REGS[4][18] , \REGS[4][17] ,
         \REGS[4][16] , \REGS[4][15] , \REGS[4][14] , \REGS[4][13] ,
         \REGS[4][12] , \REGS[4][11] , \REGS[4][10] , \REGS[4][9] ,
         \REGS[4][8] , \REGS[4][7] , \REGS[4][6] , \REGS[4][5] , \REGS[4][4] ,
         \REGS[4][3] , \REGS[4][2] , \REGS[4][1] , \REGS[4][0] , \REGS[5][31] ,
         \REGS[5][30] , \REGS[5][29] , \REGS[5][28] , \REGS[5][27] ,
         \REGS[5][26] , \REGS[5][25] , \REGS[5][24] , \REGS[5][23] ,
         \REGS[5][22] , \REGS[5][21] , \REGS[5][20] , \REGS[5][19] ,
         \REGS[5][18] , \REGS[5][17] , \REGS[5][16] , \REGS[5][15] ,
         \REGS[5][14] , \REGS[5][13] , \REGS[5][12] , \REGS[5][11] ,
         \REGS[5][10] , \REGS[5][9] , \REGS[5][8] , \REGS[5][7] , \REGS[5][6] ,
         \REGS[5][5] , \REGS[5][4] , \REGS[5][3] , \REGS[5][2] , \REGS[5][1] ,
         \REGS[5][0] , \REGS[6][31] , \REGS[6][30] , \REGS[6][29] ,
         \REGS[6][28] , \REGS[6][27] , \REGS[6][26] , \REGS[6][25] ,
         \REGS[6][24] , \REGS[6][23] , \REGS[6][22] , \REGS[6][21] ,
         \REGS[6][20] , \REGS[6][19] , \REGS[6][18] , \REGS[6][17] ,
         \REGS[6][16] , \REGS[6][15] , \REGS[6][14] , \REGS[6][13] ,
         \REGS[6][12] , \REGS[6][11] , \REGS[6][10] , \REGS[6][9] ,
         \REGS[6][8] , \REGS[6][7] , \REGS[6][6] , \REGS[6][5] , \REGS[6][4] ,
         \REGS[6][3] , \REGS[6][2] , \REGS[6][1] , \REGS[6][0] , \REGS[7][31] ,
         \REGS[7][30] , \REGS[7][29] , \REGS[7][28] , \REGS[7][27] ,
         \REGS[7][26] , \REGS[7][25] , \REGS[7][24] , \REGS[7][23] ,
         \REGS[7][22] , \REGS[7][21] , \REGS[7][20] , \REGS[7][19] ,
         \REGS[7][18] , \REGS[7][17] , \REGS[7][16] , \REGS[7][15] ,
         \REGS[7][14] , \REGS[7][13] , \REGS[7][12] , \REGS[7][11] ,
         \REGS[7][10] , \REGS[7][9] , \REGS[7][8] , \REGS[7][7] , \REGS[7][6] ,
         \REGS[7][5] , \REGS[7][4] , \REGS[7][3] , \REGS[7][2] , \REGS[7][1] ,
         \REGS[7][0] , \REGS[8][31] , \REGS[8][30] , \REGS[8][29] ,
         \REGS[8][28] , \REGS[8][27] , \REGS[8][26] , \REGS[8][25] ,
         \REGS[8][24] , \REGS[8][23] , \REGS[8][22] , \REGS[8][21] ,
         \REGS[8][20] , \REGS[8][19] , \REGS[8][18] , \REGS[8][17] ,
         \REGS[8][16] , \REGS[8][15] , \REGS[8][14] , \REGS[8][13] ,
         \REGS[8][12] , \REGS[8][11] , \REGS[8][10] , \REGS[8][9] ,
         \REGS[8][8] , \REGS[8][7] , \REGS[8][6] , \REGS[8][5] , \REGS[8][4] ,
         \REGS[8][3] , \REGS[8][2] , \REGS[8][1] , \REGS[8][0] , \REGS[9][31] ,
         \REGS[9][30] , \REGS[9][29] , \REGS[9][28] , \REGS[9][27] ,
         \REGS[9][26] , \REGS[9][25] , \REGS[9][24] , \REGS[9][23] ,
         \REGS[9][22] , \REGS[9][21] , \REGS[9][20] , \REGS[9][19] ,
         \REGS[9][18] , \REGS[9][17] , \REGS[9][16] , \REGS[9][15] ,
         \REGS[9][14] , \REGS[9][13] , \REGS[9][12] , \REGS[9][11] ,
         \REGS[9][10] , \REGS[9][9] , \REGS[9][8] , \REGS[9][7] , \REGS[9][6] ,
         \REGS[9][5] , \REGS[9][4] , \REGS[9][3] , \REGS[9][2] , \REGS[9][1] ,
         \REGS[9][0] , \REGS[10][31] , \REGS[10][30] , \REGS[10][29] ,
         \REGS[10][28] , \REGS[10][27] , \REGS[10][26] , \REGS[10][25] ,
         \REGS[10][24] , \REGS[10][23] , \REGS[10][22] , \REGS[10][21] ,
         \REGS[10][20] , \REGS[10][19] , \REGS[10][18] , \REGS[10][17] ,
         \REGS[10][16] , \REGS[10][15] , \REGS[10][14] , \REGS[10][13] ,
         \REGS[10][12] , \REGS[10][11] , \REGS[10][10] , \REGS[10][9] ,
         \REGS[10][8] , \REGS[10][7] , \REGS[10][6] , \REGS[10][5] ,
         \REGS[10][4] , \REGS[10][3] , \REGS[10][2] , \REGS[10][1] ,
         \REGS[10][0] , \REGS[11][31] , \REGS[11][30] , \REGS[11][29] ,
         \REGS[11][28] , \REGS[11][27] , \REGS[11][26] , \REGS[11][25] ,
         \REGS[11][24] , \REGS[11][23] , \REGS[11][22] , \REGS[11][21] ,
         \REGS[11][20] , \REGS[11][19] , \REGS[11][18] , \REGS[11][17] ,
         \REGS[11][16] , \REGS[11][15] , \REGS[11][14] , \REGS[11][13] ,
         \REGS[11][12] , \REGS[11][11] , \REGS[11][10] , \REGS[11][9] ,
         \REGS[11][8] , \REGS[11][7] , \REGS[11][6] , \REGS[11][5] ,
         \REGS[11][4] , \REGS[11][3] , \REGS[11][2] , \REGS[11][1] ,
         \REGS[11][0] , \REGS[12][31] , \REGS[12][30] , \REGS[12][29] ,
         \REGS[12][28] , \REGS[12][27] , \REGS[12][26] , \REGS[12][25] ,
         \REGS[12][24] , \REGS[12][23] , \REGS[12][22] , \REGS[12][21] ,
         \REGS[12][20] , \REGS[12][19] , \REGS[12][18] , \REGS[12][17] ,
         \REGS[12][16] , \REGS[12][15] , \REGS[12][14] , \REGS[12][13] ,
         \REGS[12][12] , \REGS[12][11] , \REGS[12][10] , \REGS[12][9] ,
         \REGS[12][8] , \REGS[12][7] , \REGS[12][6] , \REGS[12][5] ,
         \REGS[12][4] , \REGS[12][3] , \REGS[12][2] , \REGS[12][1] ,
         \REGS[12][0] , \REGS[13][31] , \REGS[13][30] , \REGS[13][29] ,
         \REGS[13][28] , \REGS[13][27] , \REGS[13][26] , \REGS[13][25] ,
         \REGS[13][24] , \REGS[13][23] , \REGS[13][22] , \REGS[13][21] ,
         \REGS[13][20] , \REGS[13][19] , \REGS[13][18] , \REGS[13][17] ,
         \REGS[13][16] , \REGS[13][15] , \REGS[13][14] , \REGS[13][13] ,
         \REGS[13][12] , \REGS[13][11] , \REGS[13][10] , \REGS[13][9] ,
         \REGS[13][8] , \REGS[13][7] , \REGS[13][6] , \REGS[13][5] ,
         \REGS[13][4] , \REGS[13][3] , \REGS[13][2] , \REGS[13][1] ,
         \REGS[13][0] , \REGS[14][31] , \REGS[14][30] , \REGS[14][29] ,
         \REGS[14][28] , \REGS[14][27] , \REGS[14][26] , \REGS[14][25] ,
         \REGS[14][24] , \REGS[14][23] , \REGS[14][22] , \REGS[14][21] ,
         \REGS[14][20] , \REGS[14][19] , \REGS[14][18] , \REGS[14][17] ,
         \REGS[14][16] , \REGS[14][15] , \REGS[14][14] , \REGS[14][13] ,
         \REGS[14][12] , \REGS[14][11] , \REGS[14][10] , \REGS[14][9] ,
         \REGS[14][8] , \REGS[14][7] , \REGS[14][6] , \REGS[14][5] ,
         \REGS[14][4] , \REGS[14][3] , \REGS[14][2] , \REGS[14][1] ,
         \REGS[14][0] , \REGS[15][31] , \REGS[15][30] , \REGS[15][29] ,
         \REGS[15][28] , \REGS[15][27] , \REGS[15][26] , \REGS[15][25] ,
         \REGS[15][24] , \REGS[15][23] , \REGS[15][22] , \REGS[15][21] ,
         \REGS[15][20] , \REGS[15][19] , \REGS[15][18] , \REGS[15][17] ,
         \REGS[15][16] , \REGS[15][15] , \REGS[15][14] , \REGS[15][13] ,
         \REGS[15][12] , \REGS[15][11] , \REGS[15][10] , \REGS[15][9] ,
         \REGS[15][8] , \REGS[15][7] , \REGS[15][6] , \REGS[15][5] ,
         \REGS[15][4] , \REGS[15][3] , \REGS[15][2] , \REGS[15][1] ,
         \REGS[15][0] , \REGS[16][31] , \REGS[16][30] , \REGS[16][29] ,
         \REGS[16][28] , \REGS[16][27] , \REGS[16][26] , \REGS[16][25] ,
         \REGS[16][24] , \REGS[16][23] , \REGS[16][22] , \REGS[16][21] ,
         \REGS[16][20] , \REGS[16][19] , \REGS[16][18] , \REGS[16][17] ,
         \REGS[16][16] , \REGS[16][15] , \REGS[16][14] , \REGS[16][13] ,
         \REGS[16][12] , \REGS[16][11] , \REGS[16][10] , \REGS[16][9] ,
         \REGS[16][8] , \REGS[16][7] , \REGS[16][6] , \REGS[16][5] ,
         \REGS[16][4] , \REGS[16][3] , \REGS[16][2] , \REGS[16][1] ,
         \REGS[16][0] , \REGS[17][31] , \REGS[17][30] , \REGS[17][29] ,
         \REGS[17][28] , \REGS[17][27] , \REGS[17][26] , \REGS[17][25] ,
         \REGS[17][24] , \REGS[17][23] , \REGS[17][22] , \REGS[17][21] ,
         \REGS[17][20] , \REGS[17][19] , \REGS[17][18] , \REGS[17][17] ,
         \REGS[17][16] , \REGS[17][15] , \REGS[17][14] , \REGS[17][13] ,
         \REGS[17][12] , \REGS[17][11] , \REGS[17][10] , \REGS[17][9] ,
         \REGS[17][8] , \REGS[17][7] , \REGS[17][6] , \REGS[17][5] ,
         \REGS[17][4] , \REGS[17][3] , \REGS[17][2] , \REGS[17][1] ,
         \REGS[17][0] , \REGS[18][31] , \REGS[18][30] , \REGS[18][29] ,
         \REGS[18][28] , \REGS[18][27] , \REGS[18][26] , \REGS[18][25] ,
         \REGS[18][24] , \REGS[18][23] , \REGS[18][22] , \REGS[18][21] ,
         \REGS[18][20] , \REGS[18][19] , \REGS[18][18] , \REGS[18][17] ,
         \REGS[18][16] , \REGS[18][15] , \REGS[18][14] , \REGS[18][13] ,
         \REGS[18][12] , \REGS[18][11] , \REGS[18][10] , \REGS[18][9] ,
         \REGS[18][8] , \REGS[18][7] , \REGS[18][6] , \REGS[18][5] ,
         \REGS[18][4] , \REGS[18][3] , \REGS[18][2] , \REGS[18][1] ,
         \REGS[18][0] , \REGS[19][31] , \REGS[19][30] , \REGS[19][29] ,
         \REGS[19][28] , \REGS[19][27] , \REGS[19][26] , \REGS[19][25] ,
         \REGS[19][24] , \REGS[19][23] , \REGS[19][22] , \REGS[19][21] ,
         \REGS[19][20] , \REGS[19][19] , \REGS[19][18] , \REGS[19][17] ,
         \REGS[19][16] , \REGS[19][15] , \REGS[19][14] , \REGS[19][13] ,
         \REGS[19][12] , \REGS[19][11] , \REGS[19][10] , \REGS[19][9] ,
         \REGS[19][8] , \REGS[19][7] , \REGS[19][6] , \REGS[19][5] ,
         \REGS[19][4] , \REGS[19][3] , \REGS[19][2] , \REGS[19][1] ,
         \REGS[19][0] , \REGS[20][31] , \REGS[20][30] , \REGS[20][29] ,
         \REGS[20][28] , \REGS[20][27] , \REGS[20][26] , \REGS[20][25] ,
         \REGS[20][24] , \REGS[20][23] , \REGS[20][22] , \REGS[20][21] ,
         \REGS[20][20] , \REGS[20][19] , \REGS[20][18] , \REGS[20][17] ,
         \REGS[20][16] , \REGS[20][15] , \REGS[20][14] , \REGS[20][13] ,
         \REGS[20][12] , \REGS[20][11] , \REGS[20][10] , \REGS[20][9] ,
         \REGS[20][8] , \REGS[20][7] , \REGS[20][6] , \REGS[20][5] ,
         \REGS[20][4] , \REGS[20][3] , \REGS[20][2] , \REGS[20][1] ,
         \REGS[20][0] , \REGS[21][31] , \REGS[21][30] , \REGS[21][29] ,
         \REGS[21][28] , \REGS[21][27] , \REGS[21][26] , \REGS[21][25] ,
         \REGS[21][24] , \REGS[21][23] , \REGS[21][22] , \REGS[21][21] ,
         \REGS[21][20] , \REGS[21][19] , \REGS[21][18] , \REGS[21][17] ,
         \REGS[21][16] , \REGS[21][15] , \REGS[21][14] , \REGS[21][13] ,
         \REGS[21][12] , \REGS[21][11] , \REGS[21][10] , \REGS[21][9] ,
         \REGS[21][8] , \REGS[21][7] , \REGS[21][6] , \REGS[21][5] ,
         \REGS[21][4] , \REGS[21][3] , \REGS[21][2] , \REGS[21][1] ,
         \REGS[21][0] , \REGS[22][31] , \REGS[22][30] , \REGS[22][29] ,
         \REGS[22][28] , \REGS[22][27] , \REGS[22][26] , \REGS[22][25] ,
         \REGS[22][24] , \REGS[22][23] , \REGS[22][22] , \REGS[22][21] ,
         \REGS[22][20] , \REGS[22][19] , \REGS[22][18] , \REGS[22][17] ,
         \REGS[22][16] , \REGS[22][15] , \REGS[22][14] , \REGS[22][13] ,
         \REGS[22][12] , \REGS[22][11] , \REGS[22][10] , \REGS[22][9] ,
         \REGS[22][8] , \REGS[22][7] , \REGS[22][6] , \REGS[22][5] ,
         \REGS[22][4] , \REGS[22][3] , \REGS[22][2] , \REGS[22][1] ,
         \REGS[22][0] , \REGS[23][31] , \REGS[23][30] , \REGS[23][29] ,
         \REGS[23][28] , \REGS[23][27] , \REGS[23][26] , \REGS[23][25] ,
         \REGS[23][24] , \REGS[23][23] , \REGS[23][22] , \REGS[23][21] ,
         \REGS[23][20] , \REGS[23][19] , \REGS[23][18] , \REGS[23][17] ,
         \REGS[23][16] , \REGS[23][15] , \REGS[23][14] , \REGS[23][13] ,
         \REGS[23][12] , \REGS[23][11] , \REGS[23][10] , \REGS[23][9] ,
         \REGS[23][8] , \REGS[23][7] , \REGS[23][6] , \REGS[23][5] ,
         \REGS[23][4] , \REGS[23][3] , \REGS[23][2] , \REGS[23][1] ,
         \REGS[23][0] , \REGS[24][31] , \REGS[24][30] , \REGS[24][29] ,
         \REGS[24][28] , \REGS[24][27] , \REGS[24][26] , \REGS[24][25] ,
         \REGS[24][24] , \REGS[24][23] , \REGS[24][22] , \REGS[24][21] ,
         \REGS[24][20] , \REGS[24][19] , \REGS[24][18] , \REGS[24][17] ,
         \REGS[24][16] , \REGS[24][15] , \REGS[24][14] , \REGS[24][13] ,
         \REGS[24][12] , \REGS[24][11] , \REGS[24][10] , \REGS[24][9] ,
         \REGS[24][8] , \REGS[24][7] , \REGS[24][6] , \REGS[24][5] ,
         \REGS[24][4] , \REGS[24][3] , \REGS[24][2] , \REGS[24][1] ,
         \REGS[24][0] , \REGS[25][31] , \REGS[25][30] , \REGS[25][29] ,
         \REGS[25][28] , \REGS[25][27] , \REGS[25][26] , \REGS[25][25] ,
         \REGS[25][24] , \REGS[25][23] , \REGS[25][22] , \REGS[25][21] ,
         \REGS[25][20] , \REGS[25][19] , \REGS[25][18] , \REGS[25][17] ,
         \REGS[25][16] , \REGS[25][15] , \REGS[25][14] , \REGS[25][13] ,
         \REGS[25][12] , \REGS[25][11] , \REGS[25][10] , \REGS[25][9] ,
         \REGS[25][8] , \REGS[25][7] , \REGS[25][6] , \REGS[25][5] ,
         \REGS[25][4] , \REGS[25][3] , \REGS[25][2] , \REGS[25][1] ,
         \REGS[25][0] , \REGS[26][31] , \REGS[26][30] , \REGS[26][29] ,
         \REGS[26][28] , \REGS[26][27] , \REGS[26][26] , \REGS[26][25] ,
         \REGS[26][24] , \REGS[26][23] , \REGS[26][22] , \REGS[26][21] ,
         \REGS[26][20] , \REGS[26][19] , \REGS[26][18] , \REGS[26][17] ,
         \REGS[26][16] , \REGS[26][15] , \REGS[26][14] , \REGS[26][13] ,
         \REGS[26][12] , \REGS[26][11] , \REGS[26][10] , \REGS[26][9] ,
         \REGS[26][8] , \REGS[26][7] , \REGS[26][6] , \REGS[26][5] ,
         \REGS[26][4] , \REGS[26][3] , \REGS[26][2] , \REGS[26][1] ,
         \REGS[26][0] , \REGS[27][31] , \REGS[27][30] , \REGS[27][29] ,
         \REGS[27][28] , \REGS[27][27] , \REGS[27][26] , \REGS[27][25] ,
         \REGS[27][24] , \REGS[27][23] , \REGS[27][22] , \REGS[27][21] ,
         \REGS[27][20] , \REGS[27][19] , \REGS[27][18] , \REGS[27][17] ,
         \REGS[27][16] , \REGS[27][15] , \REGS[27][14] , \REGS[27][13] ,
         \REGS[27][12] , \REGS[27][11] , \REGS[27][10] , \REGS[27][9] ,
         \REGS[27][8] , \REGS[27][7] , \REGS[27][6] , \REGS[27][5] ,
         \REGS[27][4] , \REGS[27][3] , \REGS[27][2] , \REGS[27][1] ,
         \REGS[27][0] , \REGS[28][31] , \REGS[28][30] , \REGS[28][29] ,
         \REGS[28][28] , \REGS[28][27] , \REGS[28][26] , \REGS[28][25] ,
         \REGS[28][24] , \REGS[28][23] , \REGS[28][22] , \REGS[28][21] ,
         \REGS[28][20] , \REGS[28][19] , \REGS[28][18] , \REGS[28][17] ,
         \REGS[28][16] , \REGS[28][15] , \REGS[28][14] , \REGS[28][13] ,
         \REGS[28][12] , \REGS[28][11] , \REGS[28][10] , \REGS[28][9] ,
         \REGS[28][8] , \REGS[28][7] , \REGS[28][6] , \REGS[28][5] ,
         \REGS[28][4] , \REGS[28][3] , \REGS[28][2] , \REGS[28][1] ,
         \REGS[28][0] , \REGS[29][31] , \REGS[29][30] , \REGS[29][29] ,
         \REGS[29][28] , \REGS[29][27] , \REGS[29][26] , \REGS[29][25] ,
         \REGS[29][24] , \REGS[29][23] , \REGS[29][22] , \REGS[29][21] ,
         \REGS[29][20] , \REGS[29][19] , \REGS[29][18] , \REGS[29][17] ,
         \REGS[29][16] , \REGS[29][15] , \REGS[29][14] , \REGS[29][13] ,
         \REGS[29][12] , \REGS[29][11] , \REGS[29][10] , \REGS[29][9] ,
         \REGS[29][8] , \REGS[29][7] , \REGS[29][6] , \REGS[29][5] ,
         \REGS[29][4] , \REGS[29][3] , \REGS[29][2] , \REGS[29][1] ,
         \REGS[29][0] , \REGS[30][31] , \REGS[30][30] , \REGS[30][29] ,
         \REGS[30][28] , \REGS[30][27] , \REGS[30][26] , \REGS[30][25] ,
         \REGS[30][24] , \REGS[30][23] , \REGS[30][22] , \REGS[30][21] ,
         \REGS[30][20] , \REGS[30][19] , \REGS[30][18] , \REGS[30][17] ,
         \REGS[30][16] , \REGS[30][15] , \REGS[30][14] , \REGS[30][13] ,
         \REGS[30][12] , \REGS[30][11] , \REGS[30][10] , \REGS[30][9] ,
         \REGS[30][8] , \REGS[30][7] , \REGS[30][6] , \REGS[30][5] ,
         \REGS[30][4] , \REGS[30][3] , \REGS[30][2] , \REGS[30][1] ,
         \REGS[30][0] , \REGS[31][31] , \REGS[31][30] , \REGS[31][29] ,
         \REGS[31][28] , \REGS[31][27] , \REGS[31][26] , \REGS[31][25] ,
         \REGS[31][24] , \REGS[31][23] , \REGS[31][22] , \REGS[31][21] ,
         \REGS[31][20] , \REGS[31][19] , \REGS[31][18] , \REGS[31][17] ,
         \REGS[31][16] , \REGS[31][15] , \REGS[31][14] , \REGS[31][13] ,
         \REGS[31][12] , \REGS[31][11] , \REGS[31][10] , \REGS[31][9] ,
         \REGS[31][8] , \REGS[31][7] , \REGS[31][6] , \REGS[31][5] ,
         \REGS[31][4] , \REGS[31][3] , \REGS[31][2] , \REGS[31][1] ,
         \REGS[31][0] , N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89,
         N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102,
         N103, N104, N105, N106, N107, N108, N109, N110, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N310, N343, N344, N346,
         N347, N348, N350, N351, N352, N354, N355, N356, N358, N359, N360,
         N362, N363, N364, N366, N367, N368, N370, N371, N372, N374, N375,
         N376, N378, N379, N380, N382, N384, N385, N386, N387, N388, N389,
         N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400,
         N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411,
         N412, N413, N414, N415, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248;

  DLL_X1 \REGS_reg[0][31]  ( .D(N415), .GN(n195), .Q(\REGS[0][31] ) );
  DLL_X1 \REGS_reg[0][30]  ( .D(N414), .GN(n195), .Q(\REGS[0][30] ) );
  DLL_X1 \REGS_reg[0][29]  ( .D(N413), .GN(n195), .Q(\REGS[0][29] ) );
  DLL_X1 \REGS_reg[0][28]  ( .D(N412), .GN(n195), .Q(\REGS[0][28] ) );
  DLL_X1 \REGS_reg[0][27]  ( .D(N411), .GN(n195), .Q(\REGS[0][27] ) );
  DLL_X1 \REGS_reg[0][26]  ( .D(N410), .GN(n195), .Q(\REGS[0][26] ) );
  DLL_X1 \REGS_reg[0][25]  ( .D(N409), .GN(n195), .Q(\REGS[0][25] ) );
  DLL_X1 \REGS_reg[0][24]  ( .D(N408), .GN(n195), .Q(\REGS[0][24] ) );
  DLL_X1 \REGS_reg[0][23]  ( .D(N407), .GN(n195), .Q(\REGS[0][23] ) );
  DLL_X1 \REGS_reg[0][22]  ( .D(N406), .GN(n195), .Q(\REGS[0][22] ) );
  DLL_X1 \REGS_reg[0][21]  ( .D(N405), .GN(n194), .Q(\REGS[0][21] ) );
  DLL_X1 \REGS_reg[0][20]  ( .D(N404), .GN(n194), .Q(\REGS[0][20] ) );
  DLL_X1 \REGS_reg[0][19]  ( .D(N403), .GN(n194), .Q(\REGS[0][19] ) );
  DLL_X1 \REGS_reg[0][18]  ( .D(N402), .GN(n194), .Q(\REGS[0][18] ) );
  DLL_X1 \REGS_reg[0][17]  ( .D(N401), .GN(n194), .Q(\REGS[0][17] ) );
  DLL_X1 \REGS_reg[0][16]  ( .D(N400), .GN(n194), .Q(\REGS[0][16] ) );
  DLL_X1 \REGS_reg[0][15]  ( .D(N399), .GN(n194), .Q(\REGS[0][15] ) );
  DLL_X1 \REGS_reg[0][14]  ( .D(N398), .GN(n194), .Q(\REGS[0][14] ) );
  DLL_X1 \REGS_reg[0][13]  ( .D(N397), .GN(n194), .Q(\REGS[0][13] ) );
  DLL_X1 \REGS_reg[0][12]  ( .D(N396), .GN(n194), .Q(\REGS[0][12] ) );
  DLL_X1 \REGS_reg[0][11]  ( .D(N395), .GN(n194), .Q(\REGS[0][11] ) );
  DLL_X1 \REGS_reg[0][10]  ( .D(N394), .GN(n193), .Q(\REGS[0][10] ) );
  DLL_X1 \REGS_reg[0][9]  ( .D(N393), .GN(n193), .Q(\REGS[0][9] ) );
  DLL_X1 \REGS_reg[0][8]  ( .D(N392), .GN(n193), .Q(\REGS[0][8] ) );
  DLL_X1 \REGS_reg[0][7]  ( .D(N391), .GN(n193), .Q(\REGS[0][7] ) );
  DLL_X1 \REGS_reg[0][6]  ( .D(N390), .GN(n193), .Q(\REGS[0][6] ) );
  DLL_X1 \REGS_reg[0][5]  ( .D(N389), .GN(n193), .Q(\REGS[0][5] ) );
  DLL_X1 \REGS_reg[0][4]  ( .D(N388), .GN(n193), .Q(\REGS[0][4] ) );
  DLL_X1 \REGS_reg[0][3]  ( .D(N387), .GN(n193), .Q(\REGS[0][3] ) );
  DLL_X1 \REGS_reg[0][2]  ( .D(N386), .GN(n193), .Q(\REGS[0][2] ) );
  DLL_X1 \REGS_reg[0][1]  ( .D(N385), .GN(n193), .Q(\REGS[0][1] ) );
  DLL_X1 \REGS_reg[0][0]  ( .D(N384), .GN(n193), .Q(\REGS[0][0] ) );
  DLH_X1 \REGS_reg[1][31]  ( .G(n297), .D(n1), .Q(\REGS[1][31] ) );
  DLH_X1 \REGS_reg[1][30]  ( .G(n297), .D(n4), .Q(\REGS[1][30] ) );
  DLH_X1 \REGS_reg[1][29]  ( .G(n297), .D(n7), .Q(\REGS[1][29] ) );
  DLH_X1 \REGS_reg[1][28]  ( .G(n297), .D(n10), .Q(\REGS[1][28] ) );
  DLH_X1 \REGS_reg[1][27]  ( .G(n297), .D(n13), .Q(\REGS[1][27] ) );
  DLH_X1 \REGS_reg[1][26]  ( .G(n297), .D(n16), .Q(\REGS[1][26] ) );
  DLH_X1 \REGS_reg[1][25]  ( .G(n297), .D(n19), .Q(\REGS[1][25] ) );
  DLH_X1 \REGS_reg[1][24]  ( .G(n297), .D(n22), .Q(\REGS[1][24] ) );
  DLH_X1 \REGS_reg[1][23]  ( .G(n297), .D(n25), .Q(\REGS[1][23] ) );
  DLH_X1 \REGS_reg[1][22]  ( .G(n297), .D(n28), .Q(\REGS[1][22] ) );
  DLH_X1 \REGS_reg[1][21]  ( .G(n296), .D(n31), .Q(\REGS[1][21] ) );
  DLH_X1 \REGS_reg[1][20]  ( .G(n296), .D(n34), .Q(\REGS[1][20] ) );
  DLH_X1 \REGS_reg[1][19]  ( .G(n296), .D(n37), .Q(\REGS[1][19] ) );
  DLH_X1 \REGS_reg[1][18]  ( .G(n296), .D(n40), .Q(\REGS[1][18] ) );
  DLH_X1 \REGS_reg[1][17]  ( .G(n296), .D(n43), .Q(\REGS[1][17] ) );
  DLH_X1 \REGS_reg[1][16]  ( .G(n296), .D(n46), .Q(\REGS[1][16] ) );
  DLH_X1 \REGS_reg[1][15]  ( .G(n296), .D(n49), .Q(\REGS[1][15] ) );
  DLH_X1 \REGS_reg[1][14]  ( .G(n296), .D(n52), .Q(\REGS[1][14] ) );
  DLH_X1 \REGS_reg[1][13]  ( .G(n296), .D(n55), .Q(\REGS[1][13] ) );
  DLH_X1 \REGS_reg[1][12]  ( .G(n296), .D(n58), .Q(\REGS[1][12] ) );
  DLH_X1 \REGS_reg[1][11]  ( .G(n296), .D(n61), .Q(\REGS[1][11] ) );
  DLH_X1 \REGS_reg[1][10]  ( .G(n295), .D(n64), .Q(\REGS[1][10] ) );
  DLH_X1 \REGS_reg[1][9]  ( .G(n295), .D(n67), .Q(\REGS[1][9] ) );
  DLH_X1 \REGS_reg[1][8]  ( .G(n295), .D(n70), .Q(\REGS[1][8] ) );
  DLH_X1 \REGS_reg[1][7]  ( .G(n295), .D(n73), .Q(\REGS[1][7] ) );
  DLH_X1 \REGS_reg[1][6]  ( .G(n295), .D(n76), .Q(\REGS[1][6] ) );
  DLH_X1 \REGS_reg[1][5]  ( .G(n295), .D(n79), .Q(\REGS[1][5] ) );
  DLH_X1 \REGS_reg[1][4]  ( .G(n295), .D(n82), .Q(\REGS[1][4] ) );
  DLH_X1 \REGS_reg[1][3]  ( .G(n295), .D(n85), .Q(\REGS[1][3] ) );
  DLH_X1 \REGS_reg[1][2]  ( .G(n295), .D(n88), .Q(\REGS[1][2] ) );
  DLH_X1 \REGS_reg[1][1]  ( .G(n295), .D(n91), .Q(\REGS[1][1] ) );
  DLH_X1 \REGS_reg[1][0]  ( .G(n295), .D(n94), .Q(\REGS[1][0] ) );
  DLH_X1 \REGS_reg[2][31]  ( .G(n300), .D(n1), .Q(\REGS[2][31] ) );
  DLH_X1 \REGS_reg[2][30]  ( .G(n300), .D(n4), .Q(\REGS[2][30] ) );
  DLH_X1 \REGS_reg[2][29]  ( .G(n300), .D(n7), .Q(\REGS[2][29] ) );
  DLH_X1 \REGS_reg[2][28]  ( .G(n300), .D(n10), .Q(\REGS[2][28] ) );
  DLH_X1 \REGS_reg[2][27]  ( .G(n300), .D(n13), .Q(\REGS[2][27] ) );
  DLH_X1 \REGS_reg[2][26]  ( .G(n300), .D(n16), .Q(\REGS[2][26] ) );
  DLH_X1 \REGS_reg[2][25]  ( .G(n300), .D(n19), .Q(\REGS[2][25] ) );
  DLH_X1 \REGS_reg[2][24]  ( .G(n300), .D(n22), .Q(\REGS[2][24] ) );
  DLH_X1 \REGS_reg[2][23]  ( .G(n300), .D(n25), .Q(\REGS[2][23] ) );
  DLH_X1 \REGS_reg[2][22]  ( .G(n300), .D(n28), .Q(\REGS[2][22] ) );
  DLH_X1 \REGS_reg[2][21]  ( .G(n299), .D(n31), .Q(\REGS[2][21] ) );
  DLH_X1 \REGS_reg[2][20]  ( .G(n299), .D(n34), .Q(\REGS[2][20] ) );
  DLH_X1 \REGS_reg[2][19]  ( .G(n299), .D(n37), .Q(\REGS[2][19] ) );
  DLH_X1 \REGS_reg[2][18]  ( .G(n299), .D(n40), .Q(\REGS[2][18] ) );
  DLH_X1 \REGS_reg[2][17]  ( .G(n299), .D(n43), .Q(\REGS[2][17] ) );
  DLH_X1 \REGS_reg[2][16]  ( .G(n299), .D(n46), .Q(\REGS[2][16] ) );
  DLH_X1 \REGS_reg[2][15]  ( .G(n299), .D(n49), .Q(\REGS[2][15] ) );
  DLH_X1 \REGS_reg[2][14]  ( .G(n299), .D(n52), .Q(\REGS[2][14] ) );
  DLH_X1 \REGS_reg[2][13]  ( .G(n299), .D(n55), .Q(\REGS[2][13] ) );
  DLH_X1 \REGS_reg[2][12]  ( .G(n299), .D(n58), .Q(\REGS[2][12] ) );
  DLH_X1 \REGS_reg[2][11]  ( .G(n299), .D(n61), .Q(\REGS[2][11] ) );
  DLH_X1 \REGS_reg[2][10]  ( .G(n298), .D(n64), .Q(\REGS[2][10] ) );
  DLH_X1 \REGS_reg[2][9]  ( .G(n298), .D(n67), .Q(\REGS[2][9] ) );
  DLH_X1 \REGS_reg[2][8]  ( .G(n298), .D(n70), .Q(\REGS[2][8] ) );
  DLH_X1 \REGS_reg[2][7]  ( .G(n298), .D(n73), .Q(\REGS[2][7] ) );
  DLH_X1 \REGS_reg[2][6]  ( .G(n298), .D(n76), .Q(\REGS[2][6] ) );
  DLH_X1 \REGS_reg[2][5]  ( .G(n298), .D(n79), .Q(\REGS[2][5] ) );
  DLH_X1 \REGS_reg[2][4]  ( .G(n298), .D(n82), .Q(\REGS[2][4] ) );
  DLH_X1 \REGS_reg[2][3]  ( .G(n298), .D(n85), .Q(\REGS[2][3] ) );
  DLH_X1 \REGS_reg[2][2]  ( .G(n298), .D(n88), .Q(\REGS[2][2] ) );
  DLH_X1 \REGS_reg[2][1]  ( .G(n298), .D(n91), .Q(\REGS[2][1] ) );
  DLH_X1 \REGS_reg[2][0]  ( .G(n298), .D(n94), .Q(\REGS[2][0] ) );
  DLH_X1 \REGS_reg[3][31]  ( .G(n303), .D(n1), .Q(\REGS[3][31] ) );
  DLH_X1 \REGS_reg[3][30]  ( .G(n303), .D(n4), .Q(\REGS[3][30] ) );
  DLH_X1 \REGS_reg[3][29]  ( .G(n303), .D(n7), .Q(\REGS[3][29] ) );
  DLH_X1 \REGS_reg[3][28]  ( .G(n303), .D(n10), .Q(\REGS[3][28] ) );
  DLH_X1 \REGS_reg[3][27]  ( .G(n303), .D(n13), .Q(\REGS[3][27] ) );
  DLH_X1 \REGS_reg[3][26]  ( .G(n303), .D(n16), .Q(\REGS[3][26] ) );
  DLH_X1 \REGS_reg[3][25]  ( .G(n303), .D(n19), .Q(\REGS[3][25] ) );
  DLH_X1 \REGS_reg[3][24]  ( .G(n303), .D(n22), .Q(\REGS[3][24] ) );
  DLH_X1 \REGS_reg[3][23]  ( .G(n303), .D(n25), .Q(\REGS[3][23] ) );
  DLH_X1 \REGS_reg[3][22]  ( .G(n303), .D(n28), .Q(\REGS[3][22] ) );
  DLH_X1 \REGS_reg[3][21]  ( .G(n302), .D(n31), .Q(\REGS[3][21] ) );
  DLH_X1 \REGS_reg[3][20]  ( .G(n302), .D(n34), .Q(\REGS[3][20] ) );
  DLH_X1 \REGS_reg[3][19]  ( .G(n302), .D(n37), .Q(\REGS[3][19] ) );
  DLH_X1 \REGS_reg[3][18]  ( .G(n302), .D(n40), .Q(\REGS[3][18] ) );
  DLH_X1 \REGS_reg[3][17]  ( .G(n302), .D(n43), .Q(\REGS[3][17] ) );
  DLH_X1 \REGS_reg[3][16]  ( .G(n302), .D(n46), .Q(\REGS[3][16] ) );
  DLH_X1 \REGS_reg[3][15]  ( .G(n302), .D(n49), .Q(\REGS[3][15] ) );
  DLH_X1 \REGS_reg[3][14]  ( .G(n302), .D(n52), .Q(\REGS[3][14] ) );
  DLH_X1 \REGS_reg[3][13]  ( .G(n302), .D(n55), .Q(\REGS[3][13] ) );
  DLH_X1 \REGS_reg[3][12]  ( .G(n302), .D(n58), .Q(\REGS[3][12] ) );
  DLH_X1 \REGS_reg[3][11]  ( .G(n302), .D(n61), .Q(\REGS[3][11] ) );
  DLH_X1 \REGS_reg[3][10]  ( .G(n301), .D(n64), .Q(\REGS[3][10] ) );
  DLH_X1 \REGS_reg[3][9]  ( .G(n301), .D(n67), .Q(\REGS[3][9] ) );
  DLH_X1 \REGS_reg[3][8]  ( .G(n301), .D(n70), .Q(\REGS[3][8] ) );
  DLH_X1 \REGS_reg[3][7]  ( .G(n301), .D(n73), .Q(\REGS[3][7] ) );
  DLH_X1 \REGS_reg[3][6]  ( .G(n301), .D(n76), .Q(\REGS[3][6] ) );
  DLH_X1 \REGS_reg[3][5]  ( .G(n301), .D(n79), .Q(\REGS[3][5] ) );
  DLH_X1 \REGS_reg[3][4]  ( .G(n301), .D(n82), .Q(\REGS[3][4] ) );
  DLH_X1 \REGS_reg[3][3]  ( .G(n301), .D(n85), .Q(\REGS[3][3] ) );
  DLH_X1 \REGS_reg[3][2]  ( .G(n301), .D(n88), .Q(\REGS[3][2] ) );
  DLH_X1 \REGS_reg[3][1]  ( .G(n301), .D(n91), .Q(\REGS[3][1] ) );
  DLH_X1 \REGS_reg[3][0]  ( .G(n301), .D(n94), .Q(\REGS[3][0] ) );
  DLH_X1 \REGS_reg[4][31]  ( .G(n306), .D(n1), .Q(\REGS[4][31] ) );
  DLH_X1 \REGS_reg[4][30]  ( .G(n306), .D(n4), .Q(\REGS[4][30] ) );
  DLH_X1 \REGS_reg[4][29]  ( .G(n306), .D(n7), .Q(\REGS[4][29] ) );
  DLH_X1 \REGS_reg[4][28]  ( .G(n306), .D(n10), .Q(\REGS[4][28] ) );
  DLH_X1 \REGS_reg[4][27]  ( .G(n306), .D(n13), .Q(\REGS[4][27] ) );
  DLH_X1 \REGS_reg[4][26]  ( .G(n306), .D(n16), .Q(\REGS[4][26] ) );
  DLH_X1 \REGS_reg[4][25]  ( .G(n306), .D(n19), .Q(\REGS[4][25] ) );
  DLH_X1 \REGS_reg[4][24]  ( .G(n306), .D(n22), .Q(\REGS[4][24] ) );
  DLH_X1 \REGS_reg[4][23]  ( .G(n306), .D(n25), .Q(\REGS[4][23] ) );
  DLH_X1 \REGS_reg[4][22]  ( .G(n306), .D(n28), .Q(\REGS[4][22] ) );
  DLH_X1 \REGS_reg[4][21]  ( .G(n305), .D(n31), .Q(\REGS[4][21] ) );
  DLH_X1 \REGS_reg[4][20]  ( .G(n305), .D(n34), .Q(\REGS[4][20] ) );
  DLH_X1 \REGS_reg[4][19]  ( .G(n305), .D(n37), .Q(\REGS[4][19] ) );
  DLH_X1 \REGS_reg[4][18]  ( .G(n305), .D(n40), .Q(\REGS[4][18] ) );
  DLH_X1 \REGS_reg[4][17]  ( .G(n305), .D(n43), .Q(\REGS[4][17] ) );
  DLH_X1 \REGS_reg[4][16]  ( .G(n305), .D(n46), .Q(\REGS[4][16] ) );
  DLH_X1 \REGS_reg[4][15]  ( .G(n305), .D(n49), .Q(\REGS[4][15] ) );
  DLH_X1 \REGS_reg[4][14]  ( .G(n305), .D(n52), .Q(\REGS[4][14] ) );
  DLH_X1 \REGS_reg[4][13]  ( .G(n305), .D(n55), .Q(\REGS[4][13] ) );
  DLH_X1 \REGS_reg[4][12]  ( .G(n305), .D(n58), .Q(\REGS[4][12] ) );
  DLH_X1 \REGS_reg[4][11]  ( .G(n305), .D(n61), .Q(\REGS[4][11] ) );
  DLH_X1 \REGS_reg[4][10]  ( .G(n304), .D(n64), .Q(\REGS[4][10] ) );
  DLH_X1 \REGS_reg[4][9]  ( .G(n304), .D(n67), .Q(\REGS[4][9] ) );
  DLH_X1 \REGS_reg[4][8]  ( .G(n304), .D(n70), .Q(\REGS[4][8] ) );
  DLH_X1 \REGS_reg[4][7]  ( .G(n304), .D(n73), .Q(\REGS[4][7] ) );
  DLH_X1 \REGS_reg[4][6]  ( .G(n304), .D(n76), .Q(\REGS[4][6] ) );
  DLH_X1 \REGS_reg[4][5]  ( .G(n304), .D(n79), .Q(\REGS[4][5] ) );
  DLH_X1 \REGS_reg[4][4]  ( .G(n304), .D(n82), .Q(\REGS[4][4] ) );
  DLH_X1 \REGS_reg[4][3]  ( .G(n304), .D(n85), .Q(\REGS[4][3] ) );
  DLH_X1 \REGS_reg[4][2]  ( .G(n304), .D(n88), .Q(\REGS[4][2] ) );
  DLH_X1 \REGS_reg[4][1]  ( .G(n304), .D(n91), .Q(\REGS[4][1] ) );
  DLH_X1 \REGS_reg[4][0]  ( .G(n304), .D(n94), .Q(\REGS[4][0] ) );
  DLH_X1 \REGS_reg[5][31]  ( .G(n309), .D(n1), .Q(\REGS[5][31] ) );
  DLH_X1 \REGS_reg[5][30]  ( .G(n309), .D(n4), .Q(\REGS[5][30] ) );
  DLH_X1 \REGS_reg[5][29]  ( .G(n309), .D(n7), .Q(\REGS[5][29] ) );
  DLH_X1 \REGS_reg[5][28]  ( .G(n309), .D(n10), .Q(\REGS[5][28] ) );
  DLH_X1 \REGS_reg[5][27]  ( .G(n309), .D(n13), .Q(\REGS[5][27] ) );
  DLH_X1 \REGS_reg[5][26]  ( .G(n309), .D(n16), .Q(\REGS[5][26] ) );
  DLH_X1 \REGS_reg[5][25]  ( .G(n309), .D(n19), .Q(\REGS[5][25] ) );
  DLH_X1 \REGS_reg[5][24]  ( .G(n309), .D(n22), .Q(\REGS[5][24] ) );
  DLH_X1 \REGS_reg[5][23]  ( .G(n309), .D(n25), .Q(\REGS[5][23] ) );
  DLH_X1 \REGS_reg[5][22]  ( .G(n309), .D(n28), .Q(\REGS[5][22] ) );
  DLH_X1 \REGS_reg[5][21]  ( .G(n308), .D(n31), .Q(\REGS[5][21] ) );
  DLH_X1 \REGS_reg[5][20]  ( .G(n308), .D(n34), .Q(\REGS[5][20] ) );
  DLH_X1 \REGS_reg[5][19]  ( .G(n308), .D(n37), .Q(\REGS[5][19] ) );
  DLH_X1 \REGS_reg[5][18]  ( .G(n308), .D(n40), .Q(\REGS[5][18] ) );
  DLH_X1 \REGS_reg[5][17]  ( .G(n308), .D(n43), .Q(\REGS[5][17] ) );
  DLH_X1 \REGS_reg[5][16]  ( .G(n308), .D(n46), .Q(\REGS[5][16] ) );
  DLH_X1 \REGS_reg[5][15]  ( .G(n308), .D(n49), .Q(\REGS[5][15] ) );
  DLH_X1 \REGS_reg[5][14]  ( .G(n308), .D(n52), .Q(\REGS[5][14] ) );
  DLH_X1 \REGS_reg[5][13]  ( .G(n308), .D(n55), .Q(\REGS[5][13] ) );
  DLH_X1 \REGS_reg[5][12]  ( .G(n308), .D(n58), .Q(\REGS[5][12] ) );
  DLH_X1 \REGS_reg[5][11]  ( .G(n308), .D(n61), .Q(\REGS[5][11] ) );
  DLH_X1 \REGS_reg[5][10]  ( .G(n307), .D(n64), .Q(\REGS[5][10] ) );
  DLH_X1 \REGS_reg[5][9]  ( .G(n307), .D(n67), .Q(\REGS[5][9] ) );
  DLH_X1 \REGS_reg[5][8]  ( .G(n307), .D(n70), .Q(\REGS[5][8] ) );
  DLH_X1 \REGS_reg[5][7]  ( .G(n307), .D(n73), .Q(\REGS[5][7] ) );
  DLH_X1 \REGS_reg[5][6]  ( .G(n307), .D(n76), .Q(\REGS[5][6] ) );
  DLH_X1 \REGS_reg[5][5]  ( .G(n307), .D(n79), .Q(\REGS[5][5] ) );
  DLH_X1 \REGS_reg[5][4]  ( .G(n307), .D(n82), .Q(\REGS[5][4] ) );
  DLH_X1 \REGS_reg[5][3]  ( .G(n307), .D(n85), .Q(\REGS[5][3] ) );
  DLH_X1 \REGS_reg[5][2]  ( .G(n307), .D(n88), .Q(\REGS[5][2] ) );
  DLH_X1 \REGS_reg[5][1]  ( .G(n307), .D(n91), .Q(\REGS[5][1] ) );
  DLH_X1 \REGS_reg[5][0]  ( .G(n307), .D(n94), .Q(\REGS[5][0] ) );
  DLH_X1 \REGS_reg[6][31]  ( .G(n312), .D(n1), .Q(\REGS[6][31] ) );
  DLH_X1 \REGS_reg[6][30]  ( .G(n312), .D(n4), .Q(\REGS[6][30] ) );
  DLH_X1 \REGS_reg[6][29]  ( .G(n312), .D(n7), .Q(\REGS[6][29] ) );
  DLH_X1 \REGS_reg[6][28]  ( .G(n312), .D(n10), .Q(\REGS[6][28] ) );
  DLH_X1 \REGS_reg[6][27]  ( .G(n312), .D(n13), .Q(\REGS[6][27] ) );
  DLH_X1 \REGS_reg[6][26]  ( .G(n312), .D(n16), .Q(\REGS[6][26] ) );
  DLH_X1 \REGS_reg[6][25]  ( .G(n312), .D(n19), .Q(\REGS[6][25] ) );
  DLH_X1 \REGS_reg[6][24]  ( .G(n312), .D(n22), .Q(\REGS[6][24] ) );
  DLH_X1 \REGS_reg[6][23]  ( .G(n312), .D(n25), .Q(\REGS[6][23] ) );
  DLH_X1 \REGS_reg[6][22]  ( .G(n312), .D(n28), .Q(\REGS[6][22] ) );
  DLH_X1 \REGS_reg[6][21]  ( .G(n311), .D(n31), .Q(\REGS[6][21] ) );
  DLH_X1 \REGS_reg[6][20]  ( .G(n311), .D(n34), .Q(\REGS[6][20] ) );
  DLH_X1 \REGS_reg[6][19]  ( .G(n311), .D(n37), .Q(\REGS[6][19] ) );
  DLH_X1 \REGS_reg[6][18]  ( .G(n311), .D(n40), .Q(\REGS[6][18] ) );
  DLH_X1 \REGS_reg[6][17]  ( .G(n311), .D(n43), .Q(\REGS[6][17] ) );
  DLH_X1 \REGS_reg[6][16]  ( .G(n311), .D(n46), .Q(\REGS[6][16] ) );
  DLH_X1 \REGS_reg[6][15]  ( .G(n311), .D(n49), .Q(\REGS[6][15] ) );
  DLH_X1 \REGS_reg[6][14]  ( .G(n311), .D(n52), .Q(\REGS[6][14] ) );
  DLH_X1 \REGS_reg[6][13]  ( .G(n311), .D(n55), .Q(\REGS[6][13] ) );
  DLH_X1 \REGS_reg[6][12]  ( .G(n311), .D(n58), .Q(\REGS[6][12] ) );
  DLH_X1 \REGS_reg[6][11]  ( .G(n311), .D(n61), .Q(\REGS[6][11] ) );
  DLH_X1 \REGS_reg[6][10]  ( .G(n310), .D(n64), .Q(\REGS[6][10] ) );
  DLH_X1 \REGS_reg[6][9]  ( .G(n310), .D(n67), .Q(\REGS[6][9] ) );
  DLH_X1 \REGS_reg[6][8]  ( .G(n310), .D(n70), .Q(\REGS[6][8] ) );
  DLH_X1 \REGS_reg[6][7]  ( .G(n310), .D(n73), .Q(\REGS[6][7] ) );
  DLH_X1 \REGS_reg[6][6]  ( .G(n310), .D(n76), .Q(\REGS[6][6] ) );
  DLH_X1 \REGS_reg[6][5]  ( .G(n310), .D(n79), .Q(\REGS[6][5] ) );
  DLH_X1 \REGS_reg[6][4]  ( .G(n310), .D(n82), .Q(\REGS[6][4] ) );
  DLH_X1 \REGS_reg[6][3]  ( .G(n310), .D(n85), .Q(\REGS[6][3] ) );
  DLH_X1 \REGS_reg[6][2]  ( .G(n310), .D(n88), .Q(\REGS[6][2] ) );
  DLH_X1 \REGS_reg[6][1]  ( .G(n310), .D(n91), .Q(\REGS[6][1] ) );
  DLH_X1 \REGS_reg[6][0]  ( .G(n310), .D(n94), .Q(\REGS[6][0] ) );
  DLH_X1 \REGS_reg[7][31]  ( .G(n315), .D(n1), .Q(\REGS[7][31] ) );
  DLH_X1 \REGS_reg[7][30]  ( .G(n315), .D(n4), .Q(\REGS[7][30] ) );
  DLH_X1 \REGS_reg[7][29]  ( .G(n315), .D(n7), .Q(\REGS[7][29] ) );
  DLH_X1 \REGS_reg[7][28]  ( .G(n315), .D(n10), .Q(\REGS[7][28] ) );
  DLH_X1 \REGS_reg[7][27]  ( .G(n315), .D(n13), .Q(\REGS[7][27] ) );
  DLH_X1 \REGS_reg[7][26]  ( .G(n315), .D(n16), .Q(\REGS[7][26] ) );
  DLH_X1 \REGS_reg[7][25]  ( .G(n315), .D(n19), .Q(\REGS[7][25] ) );
  DLH_X1 \REGS_reg[7][24]  ( .G(n315), .D(n22), .Q(\REGS[7][24] ) );
  DLH_X1 \REGS_reg[7][23]  ( .G(n315), .D(n25), .Q(\REGS[7][23] ) );
  DLH_X1 \REGS_reg[7][22]  ( .G(n315), .D(n28), .Q(\REGS[7][22] ) );
  DLH_X1 \REGS_reg[7][21]  ( .G(n314), .D(n31), .Q(\REGS[7][21] ) );
  DLH_X1 \REGS_reg[7][20]  ( .G(n314), .D(n34), .Q(\REGS[7][20] ) );
  DLH_X1 \REGS_reg[7][19]  ( .G(n314), .D(n37), .Q(\REGS[7][19] ) );
  DLH_X1 \REGS_reg[7][18]  ( .G(n314), .D(n40), .Q(\REGS[7][18] ) );
  DLH_X1 \REGS_reg[7][17]  ( .G(n314), .D(n43), .Q(\REGS[7][17] ) );
  DLH_X1 \REGS_reg[7][16]  ( .G(n314), .D(n46), .Q(\REGS[7][16] ) );
  DLH_X1 \REGS_reg[7][15]  ( .G(n314), .D(n49), .Q(\REGS[7][15] ) );
  DLH_X1 \REGS_reg[7][14]  ( .G(n314), .D(n52), .Q(\REGS[7][14] ) );
  DLH_X1 \REGS_reg[7][13]  ( .G(n314), .D(n55), .Q(\REGS[7][13] ) );
  DLH_X1 \REGS_reg[7][12]  ( .G(n314), .D(n58), .Q(\REGS[7][12] ) );
  DLH_X1 \REGS_reg[7][11]  ( .G(n314), .D(n61), .Q(\REGS[7][11] ) );
  DLH_X1 \REGS_reg[7][10]  ( .G(n313), .D(n64), .Q(\REGS[7][10] ) );
  DLH_X1 \REGS_reg[7][9]  ( .G(n313), .D(n67), .Q(\REGS[7][9] ) );
  DLH_X1 \REGS_reg[7][8]  ( .G(n313), .D(n70), .Q(\REGS[7][8] ) );
  DLH_X1 \REGS_reg[7][7]  ( .G(n313), .D(n73), .Q(\REGS[7][7] ) );
  DLH_X1 \REGS_reg[7][6]  ( .G(n313), .D(n76), .Q(\REGS[7][6] ) );
  DLH_X1 \REGS_reg[7][5]  ( .G(n313), .D(n79), .Q(\REGS[7][5] ) );
  DLH_X1 \REGS_reg[7][4]  ( .G(n313), .D(n82), .Q(\REGS[7][4] ) );
  DLH_X1 \REGS_reg[7][3]  ( .G(n313), .D(n85), .Q(\REGS[7][3] ) );
  DLH_X1 \REGS_reg[7][2]  ( .G(n313), .D(n88), .Q(\REGS[7][2] ) );
  DLH_X1 \REGS_reg[7][1]  ( .G(n313), .D(n91), .Q(\REGS[7][1] ) );
  DLH_X1 \REGS_reg[7][0]  ( .G(n313), .D(n94), .Q(\REGS[7][0] ) );
  DLH_X1 \REGS_reg[8][31]  ( .G(n318), .D(n1), .Q(\REGS[8][31] ) );
  DLH_X1 \REGS_reg[8][30]  ( .G(n318), .D(n4), .Q(\REGS[8][30] ) );
  DLH_X1 \REGS_reg[8][29]  ( .G(n318), .D(n7), .Q(\REGS[8][29] ) );
  DLH_X1 \REGS_reg[8][28]  ( .G(n318), .D(n10), .Q(\REGS[8][28] ) );
  DLH_X1 \REGS_reg[8][27]  ( .G(n318), .D(n13), .Q(\REGS[8][27] ) );
  DLH_X1 \REGS_reg[8][26]  ( .G(n318), .D(n16), .Q(\REGS[8][26] ) );
  DLH_X1 \REGS_reg[8][25]  ( .G(n318), .D(n19), .Q(\REGS[8][25] ) );
  DLH_X1 \REGS_reg[8][24]  ( .G(n318), .D(n22), .Q(\REGS[8][24] ) );
  DLH_X1 \REGS_reg[8][23]  ( .G(n318), .D(n25), .Q(\REGS[8][23] ) );
  DLH_X1 \REGS_reg[8][22]  ( .G(n318), .D(n28), .Q(\REGS[8][22] ) );
  DLH_X1 \REGS_reg[8][21]  ( .G(n317), .D(n31), .Q(\REGS[8][21] ) );
  DLH_X1 \REGS_reg[8][20]  ( .G(n317), .D(n34), .Q(\REGS[8][20] ) );
  DLH_X1 \REGS_reg[8][19]  ( .G(n317), .D(n37), .Q(\REGS[8][19] ) );
  DLH_X1 \REGS_reg[8][18]  ( .G(n317), .D(n40), .Q(\REGS[8][18] ) );
  DLH_X1 \REGS_reg[8][17]  ( .G(n317), .D(n43), .Q(\REGS[8][17] ) );
  DLH_X1 \REGS_reg[8][16]  ( .G(n317), .D(n46), .Q(\REGS[8][16] ) );
  DLH_X1 \REGS_reg[8][15]  ( .G(n317), .D(n49), .Q(\REGS[8][15] ) );
  DLH_X1 \REGS_reg[8][14]  ( .G(n317), .D(n52), .Q(\REGS[8][14] ) );
  DLH_X1 \REGS_reg[8][13]  ( .G(n317), .D(n55), .Q(\REGS[8][13] ) );
  DLH_X1 \REGS_reg[8][12]  ( .G(n317), .D(n58), .Q(\REGS[8][12] ) );
  DLH_X1 \REGS_reg[8][11]  ( .G(n317), .D(n61), .Q(\REGS[8][11] ) );
  DLH_X1 \REGS_reg[8][10]  ( .G(n316), .D(n64), .Q(\REGS[8][10] ) );
  DLH_X1 \REGS_reg[8][9]  ( .G(n316), .D(n67), .Q(\REGS[8][9] ) );
  DLH_X1 \REGS_reg[8][8]  ( .G(n316), .D(n70), .Q(\REGS[8][8] ) );
  DLH_X1 \REGS_reg[8][7]  ( .G(n316), .D(n73), .Q(\REGS[8][7] ) );
  DLH_X1 \REGS_reg[8][6]  ( .G(n316), .D(n76), .Q(\REGS[8][6] ) );
  DLH_X1 \REGS_reg[8][5]  ( .G(n316), .D(n79), .Q(\REGS[8][5] ) );
  DLH_X1 \REGS_reg[8][4]  ( .G(n316), .D(n82), .Q(\REGS[8][4] ) );
  DLH_X1 \REGS_reg[8][3]  ( .G(n316), .D(n85), .Q(\REGS[8][3] ) );
  DLH_X1 \REGS_reg[8][2]  ( .G(n316), .D(n88), .Q(\REGS[8][2] ) );
  DLH_X1 \REGS_reg[8][1]  ( .G(n316), .D(n91), .Q(\REGS[8][1] ) );
  DLH_X1 \REGS_reg[8][0]  ( .G(n316), .D(n94), .Q(\REGS[8][0] ) );
  DLH_X1 \REGS_reg[9][31]  ( .G(n321), .D(n1), .Q(\REGS[9][31] ) );
  DLH_X1 \REGS_reg[9][30]  ( .G(n321), .D(n4), .Q(\REGS[9][30] ) );
  DLH_X1 \REGS_reg[9][29]  ( .G(n321), .D(n7), .Q(\REGS[9][29] ) );
  DLH_X1 \REGS_reg[9][28]  ( .G(n321), .D(n10), .Q(\REGS[9][28] ) );
  DLH_X1 \REGS_reg[9][27]  ( .G(n321), .D(n13), .Q(\REGS[9][27] ) );
  DLH_X1 \REGS_reg[9][26]  ( .G(n321), .D(n16), .Q(\REGS[9][26] ) );
  DLH_X1 \REGS_reg[9][25]  ( .G(n321), .D(n19), .Q(\REGS[9][25] ) );
  DLH_X1 \REGS_reg[9][24]  ( .G(n321), .D(n22), .Q(\REGS[9][24] ) );
  DLH_X1 \REGS_reg[9][23]  ( .G(n321), .D(n25), .Q(\REGS[9][23] ) );
  DLH_X1 \REGS_reg[9][22]  ( .G(n321), .D(n28), .Q(\REGS[9][22] ) );
  DLH_X1 \REGS_reg[9][21]  ( .G(n320), .D(n31), .Q(\REGS[9][21] ) );
  DLH_X1 \REGS_reg[9][20]  ( .G(n320), .D(n34), .Q(\REGS[9][20] ) );
  DLH_X1 \REGS_reg[9][19]  ( .G(n320), .D(n37), .Q(\REGS[9][19] ) );
  DLH_X1 \REGS_reg[9][18]  ( .G(n320), .D(n40), .Q(\REGS[9][18] ) );
  DLH_X1 \REGS_reg[9][17]  ( .G(n320), .D(n43), .Q(\REGS[9][17] ) );
  DLH_X1 \REGS_reg[9][16]  ( .G(n320), .D(n46), .Q(\REGS[9][16] ) );
  DLH_X1 \REGS_reg[9][15]  ( .G(n320), .D(n49), .Q(\REGS[9][15] ) );
  DLH_X1 \REGS_reg[9][14]  ( .G(n320), .D(n52), .Q(\REGS[9][14] ) );
  DLH_X1 \REGS_reg[9][13]  ( .G(n320), .D(n55), .Q(\REGS[9][13] ) );
  DLH_X1 \REGS_reg[9][12]  ( .G(n320), .D(n58), .Q(\REGS[9][12] ) );
  DLH_X1 \REGS_reg[9][11]  ( .G(n320), .D(n61), .Q(\REGS[9][11] ) );
  DLH_X1 \REGS_reg[9][10]  ( .G(n319), .D(n64), .Q(\REGS[9][10] ) );
  DLH_X1 \REGS_reg[9][9]  ( .G(n319), .D(n67), .Q(\REGS[9][9] ) );
  DLH_X1 \REGS_reg[9][8]  ( .G(n319), .D(n70), .Q(\REGS[9][8] ) );
  DLH_X1 \REGS_reg[9][7]  ( .G(n319), .D(n73), .Q(\REGS[9][7] ) );
  DLH_X1 \REGS_reg[9][6]  ( .G(n319), .D(n76), .Q(\REGS[9][6] ) );
  DLH_X1 \REGS_reg[9][5]  ( .G(n319), .D(n79), .Q(\REGS[9][5] ) );
  DLH_X1 \REGS_reg[9][4]  ( .G(n319), .D(n82), .Q(\REGS[9][4] ) );
  DLH_X1 \REGS_reg[9][3]  ( .G(n319), .D(n85), .Q(\REGS[9][3] ) );
  DLH_X1 \REGS_reg[9][2]  ( .G(n319), .D(n88), .Q(\REGS[9][2] ) );
  DLH_X1 \REGS_reg[9][1]  ( .G(n319), .D(n91), .Q(\REGS[9][1] ) );
  DLH_X1 \REGS_reg[9][0]  ( .G(n319), .D(n94), .Q(\REGS[9][0] ) );
  DLH_X1 \REGS_reg[10][31]  ( .G(n324), .D(n1), .Q(\REGS[10][31] ) );
  DLH_X1 \REGS_reg[10][30]  ( .G(n324), .D(n4), .Q(\REGS[10][30] ) );
  DLH_X1 \REGS_reg[10][29]  ( .G(n324), .D(n7), .Q(\REGS[10][29] ) );
  DLH_X1 \REGS_reg[10][28]  ( .G(n324), .D(n10), .Q(\REGS[10][28] ) );
  DLH_X1 \REGS_reg[10][27]  ( .G(n324), .D(n13), .Q(\REGS[10][27] ) );
  DLH_X1 \REGS_reg[10][26]  ( .G(n324), .D(n16), .Q(\REGS[10][26] ) );
  DLH_X1 \REGS_reg[10][25]  ( .G(n324), .D(n19), .Q(\REGS[10][25] ) );
  DLH_X1 \REGS_reg[10][24]  ( .G(n324), .D(n22), .Q(\REGS[10][24] ) );
  DLH_X1 \REGS_reg[10][23]  ( .G(n324), .D(n25), .Q(\REGS[10][23] ) );
  DLH_X1 \REGS_reg[10][22]  ( .G(n324), .D(n28), .Q(\REGS[10][22] ) );
  DLH_X1 \REGS_reg[10][21]  ( .G(n323), .D(n31), .Q(\REGS[10][21] ) );
  DLH_X1 \REGS_reg[10][20]  ( .G(n323), .D(n34), .Q(\REGS[10][20] ) );
  DLH_X1 \REGS_reg[10][19]  ( .G(n323), .D(n37), .Q(\REGS[10][19] ) );
  DLH_X1 \REGS_reg[10][18]  ( .G(n323), .D(n40), .Q(\REGS[10][18] ) );
  DLH_X1 \REGS_reg[10][17]  ( .G(n323), .D(n43), .Q(\REGS[10][17] ) );
  DLH_X1 \REGS_reg[10][16]  ( .G(n323), .D(n46), .Q(\REGS[10][16] ) );
  DLH_X1 \REGS_reg[10][15]  ( .G(n323), .D(n49), .Q(\REGS[10][15] ) );
  DLH_X1 \REGS_reg[10][14]  ( .G(n323), .D(n52), .Q(\REGS[10][14] ) );
  DLH_X1 \REGS_reg[10][13]  ( .G(n323), .D(n55), .Q(\REGS[10][13] ) );
  DLH_X1 \REGS_reg[10][12]  ( .G(n323), .D(n58), .Q(\REGS[10][12] ) );
  DLH_X1 \REGS_reg[10][11]  ( .G(n323), .D(n61), .Q(\REGS[10][11] ) );
  DLH_X1 \REGS_reg[10][10]  ( .G(n322), .D(n64), .Q(\REGS[10][10] ) );
  DLH_X1 \REGS_reg[10][9]  ( .G(n322), .D(n67), .Q(\REGS[10][9] ) );
  DLH_X1 \REGS_reg[10][8]  ( .G(n322), .D(n70), .Q(\REGS[10][8] ) );
  DLH_X1 \REGS_reg[10][7]  ( .G(n322), .D(n73), .Q(\REGS[10][7] ) );
  DLH_X1 \REGS_reg[10][6]  ( .G(n322), .D(n76), .Q(\REGS[10][6] ) );
  DLH_X1 \REGS_reg[10][5]  ( .G(n322), .D(n79), .Q(\REGS[10][5] ) );
  DLH_X1 \REGS_reg[10][4]  ( .G(n322), .D(n82), .Q(\REGS[10][4] ) );
  DLH_X1 \REGS_reg[10][3]  ( .G(n322), .D(n85), .Q(\REGS[10][3] ) );
  DLH_X1 \REGS_reg[10][2]  ( .G(n322), .D(n88), .Q(\REGS[10][2] ) );
  DLH_X1 \REGS_reg[10][1]  ( .G(n322), .D(n91), .Q(\REGS[10][1] ) );
  DLH_X1 \REGS_reg[10][0]  ( .G(n322), .D(n94), .Q(\REGS[10][0] ) );
  DLH_X1 \REGS_reg[11][31]  ( .G(n327), .D(n1), .Q(\REGS[11][31] ) );
  DLH_X1 \REGS_reg[11][30]  ( .G(n327), .D(n4), .Q(\REGS[11][30] ) );
  DLH_X1 \REGS_reg[11][29]  ( .G(n327), .D(n7), .Q(\REGS[11][29] ) );
  DLH_X1 \REGS_reg[11][28]  ( .G(n327), .D(n10), .Q(\REGS[11][28] ) );
  DLH_X1 \REGS_reg[11][27]  ( .G(n327), .D(n13), .Q(\REGS[11][27] ) );
  DLH_X1 \REGS_reg[11][26]  ( .G(n327), .D(n16), .Q(\REGS[11][26] ) );
  DLH_X1 \REGS_reg[11][25]  ( .G(n327), .D(n19), .Q(\REGS[11][25] ) );
  DLH_X1 \REGS_reg[11][24]  ( .G(n327), .D(n22), .Q(\REGS[11][24] ) );
  DLH_X1 \REGS_reg[11][23]  ( .G(n327), .D(n25), .Q(\REGS[11][23] ) );
  DLH_X1 \REGS_reg[11][22]  ( .G(n327), .D(n28), .Q(\REGS[11][22] ) );
  DLH_X1 \REGS_reg[11][21]  ( .G(n326), .D(n31), .Q(\REGS[11][21] ) );
  DLH_X1 \REGS_reg[11][20]  ( .G(n326), .D(n34), .Q(\REGS[11][20] ) );
  DLH_X1 \REGS_reg[11][19]  ( .G(n326), .D(n37), .Q(\REGS[11][19] ) );
  DLH_X1 \REGS_reg[11][18]  ( .G(n326), .D(n40), .Q(\REGS[11][18] ) );
  DLH_X1 \REGS_reg[11][17]  ( .G(n326), .D(n43), .Q(\REGS[11][17] ) );
  DLH_X1 \REGS_reg[11][16]  ( .G(n326), .D(n46), .Q(\REGS[11][16] ) );
  DLH_X1 \REGS_reg[11][15]  ( .G(n326), .D(n49), .Q(\REGS[11][15] ) );
  DLH_X1 \REGS_reg[11][14]  ( .G(n326), .D(n52), .Q(\REGS[11][14] ) );
  DLH_X1 \REGS_reg[11][13]  ( .G(n326), .D(n55), .Q(\REGS[11][13] ) );
  DLH_X1 \REGS_reg[11][12]  ( .G(n326), .D(n58), .Q(\REGS[11][12] ) );
  DLH_X1 \REGS_reg[11][11]  ( .G(n326), .D(n61), .Q(\REGS[11][11] ) );
  DLH_X1 \REGS_reg[11][10]  ( .G(n325), .D(n64), .Q(\REGS[11][10] ) );
  DLH_X1 \REGS_reg[11][9]  ( .G(n325), .D(n67), .Q(\REGS[11][9] ) );
  DLH_X1 \REGS_reg[11][8]  ( .G(n325), .D(n70), .Q(\REGS[11][8] ) );
  DLH_X1 \REGS_reg[11][7]  ( .G(n325), .D(n73), .Q(\REGS[11][7] ) );
  DLH_X1 \REGS_reg[11][6]  ( .G(n325), .D(n76), .Q(\REGS[11][6] ) );
  DLH_X1 \REGS_reg[11][5]  ( .G(n325), .D(n79), .Q(\REGS[11][5] ) );
  DLH_X1 \REGS_reg[11][4]  ( .G(n325), .D(n82), .Q(\REGS[11][4] ) );
  DLH_X1 \REGS_reg[11][3]  ( .G(n325), .D(n85), .Q(\REGS[11][3] ) );
  DLH_X1 \REGS_reg[11][2]  ( .G(n325), .D(n88), .Q(\REGS[11][2] ) );
  DLH_X1 \REGS_reg[11][1]  ( .G(n325), .D(n91), .Q(\REGS[11][1] ) );
  DLH_X1 \REGS_reg[11][0]  ( .G(n325), .D(n94), .Q(\REGS[11][0] ) );
  DLH_X1 \REGS_reg[12][31]  ( .G(n330), .D(n2), .Q(\REGS[12][31] ) );
  DLH_X1 \REGS_reg[12][30]  ( .G(n330), .D(n5), .Q(\REGS[12][30] ) );
  DLH_X1 \REGS_reg[12][29]  ( .G(n330), .D(n8), .Q(\REGS[12][29] ) );
  DLH_X1 \REGS_reg[12][28]  ( .G(n330), .D(n11), .Q(\REGS[12][28] ) );
  DLH_X1 \REGS_reg[12][27]  ( .G(n330), .D(n14), .Q(\REGS[12][27] ) );
  DLH_X1 \REGS_reg[12][26]  ( .G(n330), .D(n17), .Q(\REGS[12][26] ) );
  DLH_X1 \REGS_reg[12][25]  ( .G(n330), .D(n20), .Q(\REGS[12][25] ) );
  DLH_X1 \REGS_reg[12][24]  ( .G(n330), .D(n23), .Q(\REGS[12][24] ) );
  DLH_X1 \REGS_reg[12][23]  ( .G(n330), .D(n26), .Q(\REGS[12][23] ) );
  DLH_X1 \REGS_reg[12][22]  ( .G(n330), .D(n29), .Q(\REGS[12][22] ) );
  DLH_X1 \REGS_reg[12][21]  ( .G(n329), .D(n32), .Q(\REGS[12][21] ) );
  DLH_X1 \REGS_reg[12][20]  ( .G(n329), .D(n35), .Q(\REGS[12][20] ) );
  DLH_X1 \REGS_reg[12][19]  ( .G(n329), .D(n38), .Q(\REGS[12][19] ) );
  DLH_X1 \REGS_reg[12][18]  ( .G(n329), .D(n41), .Q(\REGS[12][18] ) );
  DLH_X1 \REGS_reg[12][17]  ( .G(n329), .D(n44), .Q(\REGS[12][17] ) );
  DLH_X1 \REGS_reg[12][16]  ( .G(n329), .D(n47), .Q(\REGS[12][16] ) );
  DLH_X1 \REGS_reg[12][15]  ( .G(n329), .D(n50), .Q(\REGS[12][15] ) );
  DLH_X1 \REGS_reg[12][14]  ( .G(n329), .D(n53), .Q(\REGS[12][14] ) );
  DLH_X1 \REGS_reg[12][13]  ( .G(n329), .D(n56), .Q(\REGS[12][13] ) );
  DLH_X1 \REGS_reg[12][12]  ( .G(n329), .D(n59), .Q(\REGS[12][12] ) );
  DLH_X1 \REGS_reg[12][11]  ( .G(n329), .D(n62), .Q(\REGS[12][11] ) );
  DLH_X1 \REGS_reg[12][10]  ( .G(n328), .D(n65), .Q(\REGS[12][10] ) );
  DLH_X1 \REGS_reg[12][9]  ( .G(n328), .D(n68), .Q(\REGS[12][9] ) );
  DLH_X1 \REGS_reg[12][8]  ( .G(n328), .D(n71), .Q(\REGS[12][8] ) );
  DLH_X1 \REGS_reg[12][7]  ( .G(n328), .D(n74), .Q(\REGS[12][7] ) );
  DLH_X1 \REGS_reg[12][6]  ( .G(n328), .D(n77), .Q(\REGS[12][6] ) );
  DLH_X1 \REGS_reg[12][5]  ( .G(n328), .D(n80), .Q(\REGS[12][5] ) );
  DLH_X1 \REGS_reg[12][4]  ( .G(n328), .D(n83), .Q(\REGS[12][4] ) );
  DLH_X1 \REGS_reg[12][3]  ( .G(n328), .D(n86), .Q(\REGS[12][3] ) );
  DLH_X1 \REGS_reg[12][2]  ( .G(n328), .D(n89), .Q(\REGS[12][2] ) );
  DLH_X1 \REGS_reg[12][1]  ( .G(n328), .D(n92), .Q(\REGS[12][1] ) );
  DLH_X1 \REGS_reg[12][0]  ( .G(n328), .D(n95), .Q(\REGS[12][0] ) );
  DLH_X1 \REGS_reg[13][31]  ( .G(n333), .D(n2), .Q(\REGS[13][31] ) );
  DLH_X1 \REGS_reg[13][30]  ( .G(n333), .D(n5), .Q(\REGS[13][30] ) );
  DLH_X1 \REGS_reg[13][29]  ( .G(n333), .D(n8), .Q(\REGS[13][29] ) );
  DLH_X1 \REGS_reg[13][28]  ( .G(n333), .D(n11), .Q(\REGS[13][28] ) );
  DLH_X1 \REGS_reg[13][27]  ( .G(n333), .D(n14), .Q(\REGS[13][27] ) );
  DLH_X1 \REGS_reg[13][26]  ( .G(n333), .D(n17), .Q(\REGS[13][26] ) );
  DLH_X1 \REGS_reg[13][25]  ( .G(n333), .D(n20), .Q(\REGS[13][25] ) );
  DLH_X1 \REGS_reg[13][24]  ( .G(n333), .D(n23), .Q(\REGS[13][24] ) );
  DLH_X1 \REGS_reg[13][23]  ( .G(n333), .D(n26), .Q(\REGS[13][23] ) );
  DLH_X1 \REGS_reg[13][22]  ( .G(n333), .D(n29), .Q(\REGS[13][22] ) );
  DLH_X1 \REGS_reg[13][21]  ( .G(n332), .D(n32), .Q(\REGS[13][21] ) );
  DLH_X1 \REGS_reg[13][20]  ( .G(n332), .D(n35), .Q(\REGS[13][20] ) );
  DLH_X1 \REGS_reg[13][19]  ( .G(n332), .D(n38), .Q(\REGS[13][19] ) );
  DLH_X1 \REGS_reg[13][18]  ( .G(n332), .D(n41), .Q(\REGS[13][18] ) );
  DLH_X1 \REGS_reg[13][17]  ( .G(n332), .D(n44), .Q(\REGS[13][17] ) );
  DLH_X1 \REGS_reg[13][16]  ( .G(n332), .D(n47), .Q(\REGS[13][16] ) );
  DLH_X1 \REGS_reg[13][15]  ( .G(n332), .D(n50), .Q(\REGS[13][15] ) );
  DLH_X1 \REGS_reg[13][14]  ( .G(n332), .D(n53), .Q(\REGS[13][14] ) );
  DLH_X1 \REGS_reg[13][13]  ( .G(n332), .D(n56), .Q(\REGS[13][13] ) );
  DLH_X1 \REGS_reg[13][12]  ( .G(n332), .D(n59), .Q(\REGS[13][12] ) );
  DLH_X1 \REGS_reg[13][11]  ( .G(n332), .D(n62), .Q(\REGS[13][11] ) );
  DLH_X1 \REGS_reg[13][10]  ( .G(n331), .D(n65), .Q(\REGS[13][10] ) );
  DLH_X1 \REGS_reg[13][9]  ( .G(n331), .D(n68), .Q(\REGS[13][9] ) );
  DLH_X1 \REGS_reg[13][8]  ( .G(n331), .D(n71), .Q(\REGS[13][8] ) );
  DLH_X1 \REGS_reg[13][7]  ( .G(n331), .D(n74), .Q(\REGS[13][7] ) );
  DLH_X1 \REGS_reg[13][6]  ( .G(n331), .D(n77), .Q(\REGS[13][6] ) );
  DLH_X1 \REGS_reg[13][5]  ( .G(n331), .D(n80), .Q(\REGS[13][5] ) );
  DLH_X1 \REGS_reg[13][4]  ( .G(n331), .D(n83), .Q(\REGS[13][4] ) );
  DLH_X1 \REGS_reg[13][3]  ( .G(n331), .D(n86), .Q(\REGS[13][3] ) );
  DLH_X1 \REGS_reg[13][2]  ( .G(n331), .D(n89), .Q(\REGS[13][2] ) );
  DLH_X1 \REGS_reg[13][1]  ( .G(n331), .D(n92), .Q(\REGS[13][1] ) );
  DLH_X1 \REGS_reg[13][0]  ( .G(n331), .D(n95), .Q(\REGS[13][0] ) );
  DLH_X1 \REGS_reg[14][31]  ( .G(n336), .D(n2), .Q(\REGS[14][31] ) );
  DLH_X1 \REGS_reg[14][30]  ( .G(n336), .D(n5), .Q(\REGS[14][30] ) );
  DLH_X1 \REGS_reg[14][29]  ( .G(n336), .D(n8), .Q(\REGS[14][29] ) );
  DLH_X1 \REGS_reg[14][28]  ( .G(n336), .D(n11), .Q(\REGS[14][28] ) );
  DLH_X1 \REGS_reg[14][27]  ( .G(n336), .D(n14), .Q(\REGS[14][27] ) );
  DLH_X1 \REGS_reg[14][26]  ( .G(n336), .D(n17), .Q(\REGS[14][26] ) );
  DLH_X1 \REGS_reg[14][25]  ( .G(n336), .D(n20), .Q(\REGS[14][25] ) );
  DLH_X1 \REGS_reg[14][24]  ( .G(n336), .D(n23), .Q(\REGS[14][24] ) );
  DLH_X1 \REGS_reg[14][23]  ( .G(n336), .D(n26), .Q(\REGS[14][23] ) );
  DLH_X1 \REGS_reg[14][22]  ( .G(n336), .D(n29), .Q(\REGS[14][22] ) );
  DLH_X1 \REGS_reg[14][21]  ( .G(n335), .D(n32), .Q(\REGS[14][21] ) );
  DLH_X1 \REGS_reg[14][20]  ( .G(n335), .D(n35), .Q(\REGS[14][20] ) );
  DLH_X1 \REGS_reg[14][19]  ( .G(n335), .D(n38), .Q(\REGS[14][19] ) );
  DLH_X1 \REGS_reg[14][18]  ( .G(n335), .D(n41), .Q(\REGS[14][18] ) );
  DLH_X1 \REGS_reg[14][17]  ( .G(n335), .D(n44), .Q(\REGS[14][17] ) );
  DLH_X1 \REGS_reg[14][16]  ( .G(n335), .D(n47), .Q(\REGS[14][16] ) );
  DLH_X1 \REGS_reg[14][15]  ( .G(n335), .D(n50), .Q(\REGS[14][15] ) );
  DLH_X1 \REGS_reg[14][14]  ( .G(n335), .D(n53), .Q(\REGS[14][14] ) );
  DLH_X1 \REGS_reg[14][13]  ( .G(n335), .D(n56), .Q(\REGS[14][13] ) );
  DLH_X1 \REGS_reg[14][12]  ( .G(n335), .D(n59), .Q(\REGS[14][12] ) );
  DLH_X1 \REGS_reg[14][11]  ( .G(n335), .D(n62), .Q(\REGS[14][11] ) );
  DLH_X1 \REGS_reg[14][10]  ( .G(n334), .D(n65), .Q(\REGS[14][10] ) );
  DLH_X1 \REGS_reg[14][9]  ( .G(n334), .D(n68), .Q(\REGS[14][9] ) );
  DLH_X1 \REGS_reg[14][8]  ( .G(n334), .D(n71), .Q(\REGS[14][8] ) );
  DLH_X1 \REGS_reg[14][7]  ( .G(n334), .D(n74), .Q(\REGS[14][7] ) );
  DLH_X1 \REGS_reg[14][6]  ( .G(n334), .D(n77), .Q(\REGS[14][6] ) );
  DLH_X1 \REGS_reg[14][5]  ( .G(n334), .D(n80), .Q(\REGS[14][5] ) );
  DLH_X1 \REGS_reg[14][4]  ( .G(n334), .D(n83), .Q(\REGS[14][4] ) );
  DLH_X1 \REGS_reg[14][3]  ( .G(n334), .D(n86), .Q(\REGS[14][3] ) );
  DLH_X1 \REGS_reg[14][2]  ( .G(n334), .D(n89), .Q(\REGS[14][2] ) );
  DLH_X1 \REGS_reg[14][1]  ( .G(n334), .D(n92), .Q(\REGS[14][1] ) );
  DLH_X1 \REGS_reg[14][0]  ( .G(n334), .D(n95), .Q(\REGS[14][0] ) );
  DLH_X1 \REGS_reg[15][31]  ( .G(n339), .D(n2), .Q(\REGS[15][31] ) );
  DLH_X1 \REGS_reg[15][30]  ( .G(n339), .D(n5), .Q(\REGS[15][30] ) );
  DLH_X1 \REGS_reg[15][29]  ( .G(n339), .D(n8), .Q(\REGS[15][29] ) );
  DLH_X1 \REGS_reg[15][28]  ( .G(n339), .D(n11), .Q(\REGS[15][28] ) );
  DLH_X1 \REGS_reg[15][27]  ( .G(n339), .D(n14), .Q(\REGS[15][27] ) );
  DLH_X1 \REGS_reg[15][26]  ( .G(n339), .D(n17), .Q(\REGS[15][26] ) );
  DLH_X1 \REGS_reg[15][25]  ( .G(n339), .D(n20), .Q(\REGS[15][25] ) );
  DLH_X1 \REGS_reg[15][24]  ( .G(n339), .D(n23), .Q(\REGS[15][24] ) );
  DLH_X1 \REGS_reg[15][23]  ( .G(n339), .D(n26), .Q(\REGS[15][23] ) );
  DLH_X1 \REGS_reg[15][22]  ( .G(n339), .D(n29), .Q(\REGS[15][22] ) );
  DLH_X1 \REGS_reg[15][21]  ( .G(n338), .D(n32), .Q(\REGS[15][21] ) );
  DLH_X1 \REGS_reg[15][20]  ( .G(n338), .D(n35), .Q(\REGS[15][20] ) );
  DLH_X1 \REGS_reg[15][19]  ( .G(n338), .D(n38), .Q(\REGS[15][19] ) );
  DLH_X1 \REGS_reg[15][18]  ( .G(n338), .D(n41), .Q(\REGS[15][18] ) );
  DLH_X1 \REGS_reg[15][17]  ( .G(n338), .D(n44), .Q(\REGS[15][17] ) );
  DLH_X1 \REGS_reg[15][16]  ( .G(n338), .D(n47), .Q(\REGS[15][16] ) );
  DLH_X1 \REGS_reg[15][15]  ( .G(n338), .D(n50), .Q(\REGS[15][15] ) );
  DLH_X1 \REGS_reg[15][14]  ( .G(n338), .D(n53), .Q(\REGS[15][14] ) );
  DLH_X1 \REGS_reg[15][13]  ( .G(n338), .D(n56), .Q(\REGS[15][13] ) );
  DLH_X1 \REGS_reg[15][12]  ( .G(n338), .D(n59), .Q(\REGS[15][12] ) );
  DLH_X1 \REGS_reg[15][11]  ( .G(n338), .D(n62), .Q(\REGS[15][11] ) );
  DLH_X1 \REGS_reg[15][10]  ( .G(n337), .D(n65), .Q(\REGS[15][10] ) );
  DLH_X1 \REGS_reg[15][9]  ( .G(n337), .D(n68), .Q(\REGS[15][9] ) );
  DLH_X1 \REGS_reg[15][8]  ( .G(n337), .D(n71), .Q(\REGS[15][8] ) );
  DLH_X1 \REGS_reg[15][7]  ( .G(n337), .D(n74), .Q(\REGS[15][7] ) );
  DLH_X1 \REGS_reg[15][6]  ( .G(n337), .D(n77), .Q(\REGS[15][6] ) );
  DLH_X1 \REGS_reg[15][5]  ( .G(n337), .D(n80), .Q(\REGS[15][5] ) );
  DLH_X1 \REGS_reg[15][4]  ( .G(n337), .D(n83), .Q(\REGS[15][4] ) );
  DLH_X1 \REGS_reg[15][3]  ( .G(n337), .D(n86), .Q(\REGS[15][3] ) );
  DLH_X1 \REGS_reg[15][2]  ( .G(n337), .D(n89), .Q(\REGS[15][2] ) );
  DLH_X1 \REGS_reg[15][1]  ( .G(n337), .D(n92), .Q(\REGS[15][1] ) );
  DLH_X1 \REGS_reg[15][0]  ( .G(n337), .D(n95), .Q(\REGS[15][0] ) );
  DLH_X1 \REGS_reg[16][31]  ( .G(n342), .D(n2), .Q(\REGS[16][31] ) );
  DLH_X1 \REGS_reg[16][30]  ( .G(n342), .D(n5), .Q(\REGS[16][30] ) );
  DLH_X1 \REGS_reg[16][29]  ( .G(n342), .D(n8), .Q(\REGS[16][29] ) );
  DLH_X1 \REGS_reg[16][28]  ( .G(n342), .D(n11), .Q(\REGS[16][28] ) );
  DLH_X1 \REGS_reg[16][27]  ( .G(n342), .D(n14), .Q(\REGS[16][27] ) );
  DLH_X1 \REGS_reg[16][26]  ( .G(n342), .D(n17), .Q(\REGS[16][26] ) );
  DLH_X1 \REGS_reg[16][25]  ( .G(n342), .D(n20), .Q(\REGS[16][25] ) );
  DLH_X1 \REGS_reg[16][24]  ( .G(n342), .D(n23), .Q(\REGS[16][24] ) );
  DLH_X1 \REGS_reg[16][23]  ( .G(n342), .D(n26), .Q(\REGS[16][23] ) );
  DLH_X1 \REGS_reg[16][22]  ( .G(n342), .D(n29), .Q(\REGS[16][22] ) );
  DLH_X1 \REGS_reg[16][21]  ( .G(n341), .D(n32), .Q(\REGS[16][21] ) );
  DLH_X1 \REGS_reg[16][20]  ( .G(n341), .D(n35), .Q(\REGS[16][20] ) );
  DLH_X1 \REGS_reg[16][19]  ( .G(n341), .D(n38), .Q(\REGS[16][19] ) );
  DLH_X1 \REGS_reg[16][18]  ( .G(n341), .D(n41), .Q(\REGS[16][18] ) );
  DLH_X1 \REGS_reg[16][17]  ( .G(n341), .D(n44), .Q(\REGS[16][17] ) );
  DLH_X1 \REGS_reg[16][16]  ( .G(n341), .D(n47), .Q(\REGS[16][16] ) );
  DLH_X1 \REGS_reg[16][15]  ( .G(n341), .D(n50), .Q(\REGS[16][15] ) );
  DLH_X1 \REGS_reg[16][14]  ( .G(n341), .D(n53), .Q(\REGS[16][14] ) );
  DLH_X1 \REGS_reg[16][13]  ( .G(n341), .D(n56), .Q(\REGS[16][13] ) );
  DLH_X1 \REGS_reg[16][12]  ( .G(n341), .D(n59), .Q(\REGS[16][12] ) );
  DLH_X1 \REGS_reg[16][11]  ( .G(n341), .D(n62), .Q(\REGS[16][11] ) );
  DLH_X1 \REGS_reg[16][10]  ( .G(n340), .D(n65), .Q(\REGS[16][10] ) );
  DLH_X1 \REGS_reg[16][9]  ( .G(n340), .D(n68), .Q(\REGS[16][9] ) );
  DLH_X1 \REGS_reg[16][8]  ( .G(n340), .D(n71), .Q(\REGS[16][8] ) );
  DLH_X1 \REGS_reg[16][7]  ( .G(n340), .D(n74), .Q(\REGS[16][7] ) );
  DLH_X1 \REGS_reg[16][6]  ( .G(n340), .D(n77), .Q(\REGS[16][6] ) );
  DLH_X1 \REGS_reg[16][5]  ( .G(n340), .D(n80), .Q(\REGS[16][5] ) );
  DLH_X1 \REGS_reg[16][4]  ( .G(n340), .D(n83), .Q(\REGS[16][4] ) );
  DLH_X1 \REGS_reg[16][3]  ( .G(n340), .D(n86), .Q(\REGS[16][3] ) );
  DLH_X1 \REGS_reg[16][2]  ( .G(n340), .D(n89), .Q(\REGS[16][2] ) );
  DLH_X1 \REGS_reg[16][1]  ( .G(n340), .D(n92), .Q(\REGS[16][1] ) );
  DLH_X1 \REGS_reg[16][0]  ( .G(n340), .D(n95), .Q(\REGS[16][0] ) );
  DLH_X1 \REGS_reg[17][31]  ( .G(n345), .D(n2), .Q(\REGS[17][31] ) );
  DLH_X1 \REGS_reg[17][30]  ( .G(n345), .D(n5), .Q(\REGS[17][30] ) );
  DLH_X1 \REGS_reg[17][29]  ( .G(n345), .D(n8), .Q(\REGS[17][29] ) );
  DLH_X1 \REGS_reg[17][28]  ( .G(n345), .D(n11), .Q(\REGS[17][28] ) );
  DLH_X1 \REGS_reg[17][27]  ( .G(n345), .D(n14), .Q(\REGS[17][27] ) );
  DLH_X1 \REGS_reg[17][26]  ( .G(n345), .D(n17), .Q(\REGS[17][26] ) );
  DLH_X1 \REGS_reg[17][25]  ( .G(n345), .D(n20), .Q(\REGS[17][25] ) );
  DLH_X1 \REGS_reg[17][24]  ( .G(n345), .D(n23), .Q(\REGS[17][24] ) );
  DLH_X1 \REGS_reg[17][23]  ( .G(n345), .D(n26), .Q(\REGS[17][23] ) );
  DLH_X1 \REGS_reg[17][22]  ( .G(n345), .D(n29), .Q(\REGS[17][22] ) );
  DLH_X1 \REGS_reg[17][21]  ( .G(n344), .D(n32), .Q(\REGS[17][21] ) );
  DLH_X1 \REGS_reg[17][20]  ( .G(n344), .D(n35), .Q(\REGS[17][20] ) );
  DLH_X1 \REGS_reg[17][19]  ( .G(n344), .D(n38), .Q(\REGS[17][19] ) );
  DLH_X1 \REGS_reg[17][18]  ( .G(n344), .D(n41), .Q(\REGS[17][18] ) );
  DLH_X1 \REGS_reg[17][17]  ( .G(n344), .D(n44), .Q(\REGS[17][17] ) );
  DLH_X1 \REGS_reg[17][16]  ( .G(n344), .D(n47), .Q(\REGS[17][16] ) );
  DLH_X1 \REGS_reg[17][15]  ( .G(n344), .D(n50), .Q(\REGS[17][15] ) );
  DLH_X1 \REGS_reg[17][14]  ( .G(n344), .D(n53), .Q(\REGS[17][14] ) );
  DLH_X1 \REGS_reg[17][13]  ( .G(n344), .D(n56), .Q(\REGS[17][13] ) );
  DLH_X1 \REGS_reg[17][12]  ( .G(n344), .D(n59), .Q(\REGS[17][12] ) );
  DLH_X1 \REGS_reg[17][11]  ( .G(n344), .D(n62), .Q(\REGS[17][11] ) );
  DLH_X1 \REGS_reg[17][10]  ( .G(n343), .D(n65), .Q(\REGS[17][10] ) );
  DLH_X1 \REGS_reg[17][9]  ( .G(n343), .D(n68), .Q(\REGS[17][9] ) );
  DLH_X1 \REGS_reg[17][8]  ( .G(n343), .D(n71), .Q(\REGS[17][8] ) );
  DLH_X1 \REGS_reg[17][7]  ( .G(n343), .D(n74), .Q(\REGS[17][7] ) );
  DLH_X1 \REGS_reg[17][6]  ( .G(n343), .D(n77), .Q(\REGS[17][6] ) );
  DLH_X1 \REGS_reg[17][5]  ( .G(n343), .D(n80), .Q(\REGS[17][5] ) );
  DLH_X1 \REGS_reg[17][4]  ( .G(n343), .D(n83), .Q(\REGS[17][4] ) );
  DLH_X1 \REGS_reg[17][3]  ( .G(n343), .D(n86), .Q(\REGS[17][3] ) );
  DLH_X1 \REGS_reg[17][2]  ( .G(n343), .D(n89), .Q(\REGS[17][2] ) );
  DLH_X1 \REGS_reg[17][1]  ( .G(n343), .D(n92), .Q(\REGS[17][1] ) );
  DLH_X1 \REGS_reg[17][0]  ( .G(n343), .D(n95), .Q(\REGS[17][0] ) );
  DLH_X1 \REGS_reg[18][31]  ( .G(n348), .D(n2), .Q(\REGS[18][31] ) );
  DLH_X1 \REGS_reg[18][30]  ( .G(n348), .D(n5), .Q(\REGS[18][30] ) );
  DLH_X1 \REGS_reg[18][29]  ( .G(n348), .D(n8), .Q(\REGS[18][29] ) );
  DLH_X1 \REGS_reg[18][28]  ( .G(n348), .D(n11), .Q(\REGS[18][28] ) );
  DLH_X1 \REGS_reg[18][27]  ( .G(n348), .D(n14), .Q(\REGS[18][27] ) );
  DLH_X1 \REGS_reg[18][26]  ( .G(n348), .D(n17), .Q(\REGS[18][26] ) );
  DLH_X1 \REGS_reg[18][25]  ( .G(n348), .D(n20), .Q(\REGS[18][25] ) );
  DLH_X1 \REGS_reg[18][24]  ( .G(n348), .D(n23), .Q(\REGS[18][24] ) );
  DLH_X1 \REGS_reg[18][23]  ( .G(n348), .D(n26), .Q(\REGS[18][23] ) );
  DLH_X1 \REGS_reg[18][22]  ( .G(n348), .D(n29), .Q(\REGS[18][22] ) );
  DLH_X1 \REGS_reg[18][21]  ( .G(n347), .D(n32), .Q(\REGS[18][21] ) );
  DLH_X1 \REGS_reg[18][20]  ( .G(n347), .D(n35), .Q(\REGS[18][20] ) );
  DLH_X1 \REGS_reg[18][19]  ( .G(n347), .D(n38), .Q(\REGS[18][19] ) );
  DLH_X1 \REGS_reg[18][18]  ( .G(n347), .D(n41), .Q(\REGS[18][18] ) );
  DLH_X1 \REGS_reg[18][17]  ( .G(n347), .D(n44), .Q(\REGS[18][17] ) );
  DLH_X1 \REGS_reg[18][16]  ( .G(n347), .D(n47), .Q(\REGS[18][16] ) );
  DLH_X1 \REGS_reg[18][15]  ( .G(n347), .D(n50), .Q(\REGS[18][15] ) );
  DLH_X1 \REGS_reg[18][14]  ( .G(n347), .D(n53), .Q(\REGS[18][14] ) );
  DLH_X1 \REGS_reg[18][13]  ( .G(n347), .D(n56), .Q(\REGS[18][13] ) );
  DLH_X1 \REGS_reg[18][12]  ( .G(n347), .D(n59), .Q(\REGS[18][12] ) );
  DLH_X1 \REGS_reg[18][11]  ( .G(n347), .D(n62), .Q(\REGS[18][11] ) );
  DLH_X1 \REGS_reg[18][10]  ( .G(n346), .D(n65), .Q(\REGS[18][10] ) );
  DLH_X1 \REGS_reg[18][9]  ( .G(n346), .D(n68), .Q(\REGS[18][9] ) );
  DLH_X1 \REGS_reg[18][8]  ( .G(n346), .D(n71), .Q(\REGS[18][8] ) );
  DLH_X1 \REGS_reg[18][7]  ( .G(n346), .D(n74), .Q(\REGS[18][7] ) );
  DLH_X1 \REGS_reg[18][6]  ( .G(n346), .D(n77), .Q(\REGS[18][6] ) );
  DLH_X1 \REGS_reg[18][5]  ( .G(n346), .D(n80), .Q(\REGS[18][5] ) );
  DLH_X1 \REGS_reg[18][4]  ( .G(n346), .D(n83), .Q(\REGS[18][4] ) );
  DLH_X1 \REGS_reg[18][3]  ( .G(n346), .D(n86), .Q(\REGS[18][3] ) );
  DLH_X1 \REGS_reg[18][2]  ( .G(n346), .D(n89), .Q(\REGS[18][2] ) );
  DLH_X1 \REGS_reg[18][1]  ( .G(n346), .D(n92), .Q(\REGS[18][1] ) );
  DLH_X1 \REGS_reg[18][0]  ( .G(n346), .D(n95), .Q(\REGS[18][0] ) );
  DLH_X1 \REGS_reg[19][31]  ( .G(n351), .D(n2), .Q(\REGS[19][31] ) );
  DLH_X1 \REGS_reg[19][30]  ( .G(n351), .D(n5), .Q(\REGS[19][30] ) );
  DLH_X1 \REGS_reg[19][29]  ( .G(n351), .D(n8), .Q(\REGS[19][29] ) );
  DLH_X1 \REGS_reg[19][28]  ( .G(n351), .D(n11), .Q(\REGS[19][28] ) );
  DLH_X1 \REGS_reg[19][27]  ( .G(n351), .D(n14), .Q(\REGS[19][27] ) );
  DLH_X1 \REGS_reg[19][26]  ( .G(n351), .D(n17), .Q(\REGS[19][26] ) );
  DLH_X1 \REGS_reg[19][25]  ( .G(n351), .D(n20), .Q(\REGS[19][25] ) );
  DLH_X1 \REGS_reg[19][24]  ( .G(n351), .D(n23), .Q(\REGS[19][24] ) );
  DLH_X1 \REGS_reg[19][23]  ( .G(n351), .D(n26), .Q(\REGS[19][23] ) );
  DLH_X1 \REGS_reg[19][22]  ( .G(n351), .D(n29), .Q(\REGS[19][22] ) );
  DLH_X1 \REGS_reg[19][21]  ( .G(n350), .D(n32), .Q(\REGS[19][21] ) );
  DLH_X1 \REGS_reg[19][20]  ( .G(n350), .D(n35), .Q(\REGS[19][20] ) );
  DLH_X1 \REGS_reg[19][19]  ( .G(n350), .D(n38), .Q(\REGS[19][19] ) );
  DLH_X1 \REGS_reg[19][18]  ( .G(n350), .D(n41), .Q(\REGS[19][18] ) );
  DLH_X1 \REGS_reg[19][17]  ( .G(n350), .D(n44), .Q(\REGS[19][17] ) );
  DLH_X1 \REGS_reg[19][16]  ( .G(n350), .D(n47), .Q(\REGS[19][16] ) );
  DLH_X1 \REGS_reg[19][15]  ( .G(n350), .D(n50), .Q(\REGS[19][15] ) );
  DLH_X1 \REGS_reg[19][14]  ( .G(n350), .D(n53), .Q(\REGS[19][14] ) );
  DLH_X1 \REGS_reg[19][13]  ( .G(n350), .D(n56), .Q(\REGS[19][13] ) );
  DLH_X1 \REGS_reg[19][12]  ( .G(n350), .D(n59), .Q(\REGS[19][12] ) );
  DLH_X1 \REGS_reg[19][11]  ( .G(n350), .D(n62), .Q(\REGS[19][11] ) );
  DLH_X1 \REGS_reg[19][10]  ( .G(n349), .D(n65), .Q(\REGS[19][10] ) );
  DLH_X1 \REGS_reg[19][9]  ( .G(n349), .D(n68), .Q(\REGS[19][9] ) );
  DLH_X1 \REGS_reg[19][8]  ( .G(n349), .D(n71), .Q(\REGS[19][8] ) );
  DLH_X1 \REGS_reg[19][7]  ( .G(n349), .D(n74), .Q(\REGS[19][7] ) );
  DLH_X1 \REGS_reg[19][6]  ( .G(n349), .D(n77), .Q(\REGS[19][6] ) );
  DLH_X1 \REGS_reg[19][5]  ( .G(n349), .D(n80), .Q(\REGS[19][5] ) );
  DLH_X1 \REGS_reg[19][4]  ( .G(n349), .D(n83), .Q(\REGS[19][4] ) );
  DLH_X1 \REGS_reg[19][3]  ( .G(n349), .D(n86), .Q(\REGS[19][3] ) );
  DLH_X1 \REGS_reg[19][2]  ( .G(n349), .D(n89), .Q(\REGS[19][2] ) );
  DLH_X1 \REGS_reg[19][1]  ( .G(n349), .D(n92), .Q(\REGS[19][1] ) );
  DLH_X1 \REGS_reg[19][0]  ( .G(n349), .D(n95), .Q(\REGS[19][0] ) );
  DLH_X1 \REGS_reg[20][31]  ( .G(n354), .D(n2), .Q(\REGS[20][31] ) );
  DLH_X1 \REGS_reg[20][30]  ( .G(n354), .D(n5), .Q(\REGS[20][30] ) );
  DLH_X1 \REGS_reg[20][29]  ( .G(n354), .D(n8), .Q(\REGS[20][29] ) );
  DLH_X1 \REGS_reg[20][28]  ( .G(n354), .D(n11), .Q(\REGS[20][28] ) );
  DLH_X1 \REGS_reg[20][27]  ( .G(n354), .D(n14), .Q(\REGS[20][27] ) );
  DLH_X1 \REGS_reg[20][26]  ( .G(n354), .D(n17), .Q(\REGS[20][26] ) );
  DLH_X1 \REGS_reg[20][25]  ( .G(n354), .D(n20), .Q(\REGS[20][25] ) );
  DLH_X1 \REGS_reg[20][24]  ( .G(n354), .D(n23), .Q(\REGS[20][24] ) );
  DLH_X1 \REGS_reg[20][23]  ( .G(n354), .D(n26), .Q(\REGS[20][23] ) );
  DLH_X1 \REGS_reg[20][22]  ( .G(n354), .D(n29), .Q(\REGS[20][22] ) );
  DLH_X1 \REGS_reg[20][21]  ( .G(n353), .D(n32), .Q(\REGS[20][21] ) );
  DLH_X1 \REGS_reg[20][20]  ( .G(n353), .D(n35), .Q(\REGS[20][20] ) );
  DLH_X1 \REGS_reg[20][19]  ( .G(n353), .D(n38), .Q(\REGS[20][19] ) );
  DLH_X1 \REGS_reg[20][18]  ( .G(n353), .D(n41), .Q(\REGS[20][18] ) );
  DLH_X1 \REGS_reg[20][17]  ( .G(n353), .D(n44), .Q(\REGS[20][17] ) );
  DLH_X1 \REGS_reg[20][16]  ( .G(n353), .D(n47), .Q(\REGS[20][16] ) );
  DLH_X1 \REGS_reg[20][15]  ( .G(n353), .D(n50), .Q(\REGS[20][15] ) );
  DLH_X1 \REGS_reg[20][14]  ( .G(n353), .D(n53), .Q(\REGS[20][14] ) );
  DLH_X1 \REGS_reg[20][13]  ( .G(n353), .D(n56), .Q(\REGS[20][13] ) );
  DLH_X1 \REGS_reg[20][12]  ( .G(n353), .D(n59), .Q(\REGS[20][12] ) );
  DLH_X1 \REGS_reg[20][11]  ( .G(n353), .D(n62), .Q(\REGS[20][11] ) );
  DLH_X1 \REGS_reg[20][10]  ( .G(n352), .D(n65), .Q(\REGS[20][10] ) );
  DLH_X1 \REGS_reg[20][9]  ( .G(n352), .D(n68), .Q(\REGS[20][9] ) );
  DLH_X1 \REGS_reg[20][8]  ( .G(n352), .D(n71), .Q(\REGS[20][8] ) );
  DLH_X1 \REGS_reg[20][7]  ( .G(n352), .D(n74), .Q(\REGS[20][7] ) );
  DLH_X1 \REGS_reg[20][6]  ( .G(n352), .D(n77), .Q(\REGS[20][6] ) );
  DLH_X1 \REGS_reg[20][5]  ( .G(n352), .D(n80), .Q(\REGS[20][5] ) );
  DLH_X1 \REGS_reg[20][4]  ( .G(n352), .D(n83), .Q(\REGS[20][4] ) );
  DLH_X1 \REGS_reg[20][3]  ( .G(n352), .D(n86), .Q(\REGS[20][3] ) );
  DLH_X1 \REGS_reg[20][2]  ( .G(n352), .D(n89), .Q(\REGS[20][2] ) );
  DLH_X1 \REGS_reg[20][1]  ( .G(n352), .D(n92), .Q(\REGS[20][1] ) );
  DLH_X1 \REGS_reg[20][0]  ( .G(n352), .D(n95), .Q(\REGS[20][0] ) );
  DLH_X1 \REGS_reg[21][31]  ( .G(n357), .D(n2), .Q(\REGS[21][31] ) );
  DLH_X1 \REGS_reg[21][30]  ( .G(n357), .D(n5), .Q(\REGS[21][30] ) );
  DLH_X1 \REGS_reg[21][29]  ( .G(n357), .D(n8), .Q(\REGS[21][29] ) );
  DLH_X1 \REGS_reg[21][28]  ( .G(n357), .D(n11), .Q(\REGS[21][28] ) );
  DLH_X1 \REGS_reg[21][27]  ( .G(n357), .D(n14), .Q(\REGS[21][27] ) );
  DLH_X1 \REGS_reg[21][26]  ( .G(n357), .D(n17), .Q(\REGS[21][26] ) );
  DLH_X1 \REGS_reg[21][25]  ( .G(n357), .D(n20), .Q(\REGS[21][25] ) );
  DLH_X1 \REGS_reg[21][24]  ( .G(n357), .D(n23), .Q(\REGS[21][24] ) );
  DLH_X1 \REGS_reg[21][23]  ( .G(n357), .D(n26), .Q(\REGS[21][23] ) );
  DLH_X1 \REGS_reg[21][22]  ( .G(n357), .D(n29), .Q(\REGS[21][22] ) );
  DLH_X1 \REGS_reg[21][21]  ( .G(n356), .D(n32), .Q(\REGS[21][21] ) );
  DLH_X1 \REGS_reg[21][20]  ( .G(n356), .D(n35), .Q(\REGS[21][20] ) );
  DLH_X1 \REGS_reg[21][19]  ( .G(n356), .D(n38), .Q(\REGS[21][19] ) );
  DLH_X1 \REGS_reg[21][18]  ( .G(n356), .D(n41), .Q(\REGS[21][18] ) );
  DLH_X1 \REGS_reg[21][17]  ( .G(n356), .D(n44), .Q(\REGS[21][17] ) );
  DLH_X1 \REGS_reg[21][16]  ( .G(n356), .D(n47), .Q(\REGS[21][16] ) );
  DLH_X1 \REGS_reg[21][15]  ( .G(n356), .D(n50), .Q(\REGS[21][15] ) );
  DLH_X1 \REGS_reg[21][14]  ( .G(n356), .D(n53), .Q(\REGS[21][14] ) );
  DLH_X1 \REGS_reg[21][13]  ( .G(n356), .D(n56), .Q(\REGS[21][13] ) );
  DLH_X1 \REGS_reg[21][12]  ( .G(n356), .D(n59), .Q(\REGS[21][12] ) );
  DLH_X1 \REGS_reg[21][11]  ( .G(n356), .D(n62), .Q(\REGS[21][11] ) );
  DLH_X1 \REGS_reg[21][10]  ( .G(n355), .D(n65), .Q(\REGS[21][10] ) );
  DLH_X1 \REGS_reg[21][9]  ( .G(n355), .D(n68), .Q(\REGS[21][9] ) );
  DLH_X1 \REGS_reg[21][8]  ( .G(n355), .D(n71), .Q(\REGS[21][8] ) );
  DLH_X1 \REGS_reg[21][7]  ( .G(n355), .D(n74), .Q(\REGS[21][7] ) );
  DLH_X1 \REGS_reg[21][6]  ( .G(n355), .D(n77), .Q(\REGS[21][6] ) );
  DLH_X1 \REGS_reg[21][5]  ( .G(n355), .D(n80), .Q(\REGS[21][5] ) );
  DLH_X1 \REGS_reg[21][4]  ( .G(n355), .D(n83), .Q(\REGS[21][4] ) );
  DLH_X1 \REGS_reg[21][3]  ( .G(n355), .D(n86), .Q(\REGS[21][3] ) );
  DLH_X1 \REGS_reg[21][2]  ( .G(n355), .D(n89), .Q(\REGS[21][2] ) );
  DLH_X1 \REGS_reg[21][1]  ( .G(n355), .D(n92), .Q(\REGS[21][1] ) );
  DLH_X1 \REGS_reg[21][0]  ( .G(n355), .D(n95), .Q(\REGS[21][0] ) );
  DLH_X1 \REGS_reg[22][31]  ( .G(n360), .D(n2), .Q(\REGS[22][31] ) );
  DLH_X1 \REGS_reg[22][30]  ( .G(n360), .D(n5), .Q(\REGS[22][30] ) );
  DLH_X1 \REGS_reg[22][29]  ( .G(n360), .D(n8), .Q(\REGS[22][29] ) );
  DLH_X1 \REGS_reg[22][28]  ( .G(n360), .D(n11), .Q(\REGS[22][28] ) );
  DLH_X1 \REGS_reg[22][27]  ( .G(n360), .D(n14), .Q(\REGS[22][27] ) );
  DLH_X1 \REGS_reg[22][26]  ( .G(n360), .D(n17), .Q(\REGS[22][26] ) );
  DLH_X1 \REGS_reg[22][25]  ( .G(n360), .D(n20), .Q(\REGS[22][25] ) );
  DLH_X1 \REGS_reg[22][24]  ( .G(n360), .D(n23), .Q(\REGS[22][24] ) );
  DLH_X1 \REGS_reg[22][23]  ( .G(n360), .D(n26), .Q(\REGS[22][23] ) );
  DLH_X1 \REGS_reg[22][22]  ( .G(n360), .D(n29), .Q(\REGS[22][22] ) );
  DLH_X1 \REGS_reg[22][21]  ( .G(n359), .D(n32), .Q(\REGS[22][21] ) );
  DLH_X1 \REGS_reg[22][20]  ( .G(n359), .D(n35), .Q(\REGS[22][20] ) );
  DLH_X1 \REGS_reg[22][19]  ( .G(n359), .D(n38), .Q(\REGS[22][19] ) );
  DLH_X1 \REGS_reg[22][18]  ( .G(n359), .D(n41), .Q(\REGS[22][18] ) );
  DLH_X1 \REGS_reg[22][17]  ( .G(n359), .D(n44), .Q(\REGS[22][17] ) );
  DLH_X1 \REGS_reg[22][16]  ( .G(n359), .D(n47), .Q(\REGS[22][16] ) );
  DLH_X1 \REGS_reg[22][15]  ( .G(n359), .D(n50), .Q(\REGS[22][15] ) );
  DLH_X1 \REGS_reg[22][14]  ( .G(n359), .D(n53), .Q(\REGS[22][14] ) );
  DLH_X1 \REGS_reg[22][13]  ( .G(n359), .D(n56), .Q(\REGS[22][13] ) );
  DLH_X1 \REGS_reg[22][12]  ( .G(n359), .D(n59), .Q(\REGS[22][12] ) );
  DLH_X1 \REGS_reg[22][11]  ( .G(n359), .D(n62), .Q(\REGS[22][11] ) );
  DLH_X1 \REGS_reg[22][10]  ( .G(n358), .D(n65), .Q(\REGS[22][10] ) );
  DLH_X1 \REGS_reg[22][9]  ( .G(n358), .D(n68), .Q(\REGS[22][9] ) );
  DLH_X1 \REGS_reg[22][8]  ( .G(n358), .D(n71), .Q(\REGS[22][8] ) );
  DLH_X1 \REGS_reg[22][7]  ( .G(n358), .D(n74), .Q(\REGS[22][7] ) );
  DLH_X1 \REGS_reg[22][6]  ( .G(n358), .D(n77), .Q(\REGS[22][6] ) );
  DLH_X1 \REGS_reg[22][5]  ( .G(n358), .D(n80), .Q(\REGS[22][5] ) );
  DLH_X1 \REGS_reg[22][4]  ( .G(n358), .D(n83), .Q(\REGS[22][4] ) );
  DLH_X1 \REGS_reg[22][3]  ( .G(n358), .D(n86), .Q(\REGS[22][3] ) );
  DLH_X1 \REGS_reg[22][2]  ( .G(n358), .D(n89), .Q(\REGS[22][2] ) );
  DLH_X1 \REGS_reg[22][1]  ( .G(n358), .D(n92), .Q(\REGS[22][1] ) );
  DLH_X1 \REGS_reg[22][0]  ( .G(n358), .D(n95), .Q(\REGS[22][0] ) );
  DLH_X1 \REGS_reg[23][31]  ( .G(n363), .D(n3), .Q(\REGS[23][31] ) );
  DLH_X1 \REGS_reg[23][30]  ( .G(n363), .D(n6), .Q(\REGS[23][30] ) );
  DLH_X1 \REGS_reg[23][29]  ( .G(n363), .D(n9), .Q(\REGS[23][29] ) );
  DLH_X1 \REGS_reg[23][28]  ( .G(n363), .D(n12), .Q(\REGS[23][28] ) );
  DLH_X1 \REGS_reg[23][27]  ( .G(n363), .D(n15), .Q(\REGS[23][27] ) );
  DLH_X1 \REGS_reg[23][26]  ( .G(n363), .D(n18), .Q(\REGS[23][26] ) );
  DLH_X1 \REGS_reg[23][25]  ( .G(n363), .D(n21), .Q(\REGS[23][25] ) );
  DLH_X1 \REGS_reg[23][24]  ( .G(n363), .D(n24), .Q(\REGS[23][24] ) );
  DLH_X1 \REGS_reg[23][23]  ( .G(n363), .D(n27), .Q(\REGS[23][23] ) );
  DLH_X1 \REGS_reg[23][22]  ( .G(n363), .D(n30), .Q(\REGS[23][22] ) );
  DLH_X1 \REGS_reg[23][21]  ( .G(n362), .D(n33), .Q(\REGS[23][21] ) );
  DLH_X1 \REGS_reg[23][20]  ( .G(n362), .D(n36), .Q(\REGS[23][20] ) );
  DLH_X1 \REGS_reg[23][19]  ( .G(n362), .D(n39), .Q(\REGS[23][19] ) );
  DLH_X1 \REGS_reg[23][18]  ( .G(n362), .D(n42), .Q(\REGS[23][18] ) );
  DLH_X1 \REGS_reg[23][17]  ( .G(n362), .D(n45), .Q(\REGS[23][17] ) );
  DLH_X1 \REGS_reg[23][16]  ( .G(n362), .D(n48), .Q(\REGS[23][16] ) );
  DLH_X1 \REGS_reg[23][15]  ( .G(n362), .D(n51), .Q(\REGS[23][15] ) );
  DLH_X1 \REGS_reg[23][14]  ( .G(n362), .D(n54), .Q(\REGS[23][14] ) );
  DLH_X1 \REGS_reg[23][13]  ( .G(n362), .D(n57), .Q(\REGS[23][13] ) );
  DLH_X1 \REGS_reg[23][12]  ( .G(n362), .D(n60), .Q(\REGS[23][12] ) );
  DLH_X1 \REGS_reg[23][11]  ( .G(n362), .D(n63), .Q(\REGS[23][11] ) );
  DLH_X1 \REGS_reg[23][10]  ( .G(n361), .D(n66), .Q(\REGS[23][10] ) );
  DLH_X1 \REGS_reg[23][9]  ( .G(n361), .D(n69), .Q(\REGS[23][9] ) );
  DLH_X1 \REGS_reg[23][8]  ( .G(n361), .D(n72), .Q(\REGS[23][8] ) );
  DLH_X1 \REGS_reg[23][7]  ( .G(n361), .D(n75), .Q(\REGS[23][7] ) );
  DLH_X1 \REGS_reg[23][6]  ( .G(n361), .D(n78), .Q(\REGS[23][6] ) );
  DLH_X1 \REGS_reg[23][5]  ( .G(n361), .D(n81), .Q(\REGS[23][5] ) );
  DLH_X1 \REGS_reg[23][4]  ( .G(n361), .D(n84), .Q(\REGS[23][4] ) );
  DLH_X1 \REGS_reg[23][3]  ( .G(n361), .D(n87), .Q(\REGS[23][3] ) );
  DLH_X1 \REGS_reg[23][2]  ( .G(n361), .D(n90), .Q(\REGS[23][2] ) );
  DLH_X1 \REGS_reg[23][1]  ( .G(n361), .D(n93), .Q(\REGS[23][1] ) );
  DLH_X1 \REGS_reg[23][0]  ( .G(n361), .D(n96), .Q(\REGS[23][0] ) );
  DLH_X1 \REGS_reg[24][31]  ( .G(n366), .D(n3), .Q(\REGS[24][31] ) );
  DLH_X1 \REGS_reg[24][30]  ( .G(n366), .D(n6), .Q(\REGS[24][30] ) );
  DLH_X1 \REGS_reg[24][29]  ( .G(n366), .D(n9), .Q(\REGS[24][29] ) );
  DLH_X1 \REGS_reg[24][28]  ( .G(n366), .D(n12), .Q(\REGS[24][28] ) );
  DLH_X1 \REGS_reg[24][27]  ( .G(n366), .D(n15), .Q(\REGS[24][27] ) );
  DLH_X1 \REGS_reg[24][26]  ( .G(n366), .D(n18), .Q(\REGS[24][26] ) );
  DLH_X1 \REGS_reg[24][25]  ( .G(n366), .D(n21), .Q(\REGS[24][25] ) );
  DLH_X1 \REGS_reg[24][24]  ( .G(n366), .D(n24), .Q(\REGS[24][24] ) );
  DLH_X1 \REGS_reg[24][23]  ( .G(n366), .D(n27), .Q(\REGS[24][23] ) );
  DLH_X1 \REGS_reg[24][22]  ( .G(n366), .D(n30), .Q(\REGS[24][22] ) );
  DLH_X1 \REGS_reg[24][21]  ( .G(n365), .D(n33), .Q(\REGS[24][21] ) );
  DLH_X1 \REGS_reg[24][20]  ( .G(n365), .D(n36), .Q(\REGS[24][20] ) );
  DLH_X1 \REGS_reg[24][19]  ( .G(n365), .D(n39), .Q(\REGS[24][19] ) );
  DLH_X1 \REGS_reg[24][18]  ( .G(n365), .D(n42), .Q(\REGS[24][18] ) );
  DLH_X1 \REGS_reg[24][17]  ( .G(n365), .D(n45), .Q(\REGS[24][17] ) );
  DLH_X1 \REGS_reg[24][16]  ( .G(n365), .D(n48), .Q(\REGS[24][16] ) );
  DLH_X1 \REGS_reg[24][15]  ( .G(n365), .D(n51), .Q(\REGS[24][15] ) );
  DLH_X1 \REGS_reg[24][14]  ( .G(n365), .D(n54), .Q(\REGS[24][14] ) );
  DLH_X1 \REGS_reg[24][13]  ( .G(n365), .D(n57), .Q(\REGS[24][13] ) );
  DLH_X1 \REGS_reg[24][12]  ( .G(n365), .D(n60), .Q(\REGS[24][12] ) );
  DLH_X1 \REGS_reg[24][11]  ( .G(n365), .D(n63), .Q(\REGS[24][11] ) );
  DLH_X1 \REGS_reg[24][10]  ( .G(n364), .D(n66), .Q(\REGS[24][10] ) );
  DLH_X1 \REGS_reg[24][9]  ( .G(n364), .D(n69), .Q(\REGS[24][9] ) );
  DLH_X1 \REGS_reg[24][8]  ( .G(n364), .D(n72), .Q(\REGS[24][8] ) );
  DLH_X1 \REGS_reg[24][7]  ( .G(n364), .D(n75), .Q(\REGS[24][7] ) );
  DLH_X1 \REGS_reg[24][6]  ( .G(n364), .D(n78), .Q(\REGS[24][6] ) );
  DLH_X1 \REGS_reg[24][5]  ( .G(n364), .D(n81), .Q(\REGS[24][5] ) );
  DLH_X1 \REGS_reg[24][4]  ( .G(n364), .D(n84), .Q(\REGS[24][4] ) );
  DLH_X1 \REGS_reg[24][3]  ( .G(n364), .D(n87), .Q(\REGS[24][3] ) );
  DLH_X1 \REGS_reg[24][2]  ( .G(n364), .D(n90), .Q(\REGS[24][2] ) );
  DLH_X1 \REGS_reg[24][1]  ( .G(n364), .D(n93), .Q(\REGS[24][1] ) );
  DLH_X1 \REGS_reg[24][0]  ( .G(n364), .D(n96), .Q(\REGS[24][0] ) );
  DLH_X1 \REGS_reg[25][31]  ( .G(n369), .D(n3), .Q(\REGS[25][31] ) );
  DLH_X1 \REGS_reg[25][30]  ( .G(n369), .D(n6), .Q(\REGS[25][30] ) );
  DLH_X1 \REGS_reg[25][29]  ( .G(n369), .D(n9), .Q(\REGS[25][29] ) );
  DLH_X1 \REGS_reg[25][28]  ( .G(n369), .D(n12), .Q(\REGS[25][28] ) );
  DLH_X1 \REGS_reg[25][27]  ( .G(n369), .D(n15), .Q(\REGS[25][27] ) );
  DLH_X1 \REGS_reg[25][26]  ( .G(n369), .D(n18), .Q(\REGS[25][26] ) );
  DLH_X1 \REGS_reg[25][25]  ( .G(n369), .D(n21), .Q(\REGS[25][25] ) );
  DLH_X1 \REGS_reg[25][24]  ( .G(n369), .D(n24), .Q(\REGS[25][24] ) );
  DLH_X1 \REGS_reg[25][23]  ( .G(n369), .D(n27), .Q(\REGS[25][23] ) );
  DLH_X1 \REGS_reg[25][22]  ( .G(n369), .D(n30), .Q(\REGS[25][22] ) );
  DLH_X1 \REGS_reg[25][21]  ( .G(n368), .D(n33), .Q(\REGS[25][21] ) );
  DLH_X1 \REGS_reg[25][20]  ( .G(n368), .D(n36), .Q(\REGS[25][20] ) );
  DLH_X1 \REGS_reg[25][19]  ( .G(n368), .D(n39), .Q(\REGS[25][19] ) );
  DLH_X1 \REGS_reg[25][18]  ( .G(n368), .D(n42), .Q(\REGS[25][18] ) );
  DLH_X1 \REGS_reg[25][17]  ( .G(n368), .D(n45), .Q(\REGS[25][17] ) );
  DLH_X1 \REGS_reg[25][16]  ( .G(n368), .D(n48), .Q(\REGS[25][16] ) );
  DLH_X1 \REGS_reg[25][15]  ( .G(n368), .D(n51), .Q(\REGS[25][15] ) );
  DLH_X1 \REGS_reg[25][14]  ( .G(n368), .D(n54), .Q(\REGS[25][14] ) );
  DLH_X1 \REGS_reg[25][13]  ( .G(n368), .D(n57), .Q(\REGS[25][13] ) );
  DLH_X1 \REGS_reg[25][12]  ( .G(n368), .D(n60), .Q(\REGS[25][12] ) );
  DLH_X1 \REGS_reg[25][11]  ( .G(n368), .D(n63), .Q(\REGS[25][11] ) );
  DLH_X1 \REGS_reg[25][10]  ( .G(n367), .D(n66), .Q(\REGS[25][10] ) );
  DLH_X1 \REGS_reg[25][9]  ( .G(n367), .D(n69), .Q(\REGS[25][9] ) );
  DLH_X1 \REGS_reg[25][8]  ( .G(n367), .D(n72), .Q(\REGS[25][8] ) );
  DLH_X1 \REGS_reg[25][7]  ( .G(n367), .D(n75), .Q(\REGS[25][7] ) );
  DLH_X1 \REGS_reg[25][6]  ( .G(n367), .D(n78), .Q(\REGS[25][6] ) );
  DLH_X1 \REGS_reg[25][5]  ( .G(n367), .D(n81), .Q(\REGS[25][5] ) );
  DLH_X1 \REGS_reg[25][4]  ( .G(n367), .D(n84), .Q(\REGS[25][4] ) );
  DLH_X1 \REGS_reg[25][3]  ( .G(n367), .D(n87), .Q(\REGS[25][3] ) );
  DLH_X1 \REGS_reg[25][2]  ( .G(n367), .D(n90), .Q(\REGS[25][2] ) );
  DLH_X1 \REGS_reg[25][1]  ( .G(n367), .D(n93), .Q(\REGS[25][1] ) );
  DLH_X1 \REGS_reg[25][0]  ( .G(n367), .D(n96), .Q(\REGS[25][0] ) );
  DLH_X1 \REGS_reg[26][31]  ( .G(n372), .D(n3), .Q(\REGS[26][31] ) );
  DLH_X1 \REGS_reg[26][30]  ( .G(n372), .D(n6), .Q(\REGS[26][30] ) );
  DLH_X1 \REGS_reg[26][29]  ( .G(n372), .D(n9), .Q(\REGS[26][29] ) );
  DLH_X1 \REGS_reg[26][28]  ( .G(n372), .D(n12), .Q(\REGS[26][28] ) );
  DLH_X1 \REGS_reg[26][27]  ( .G(n372), .D(n15), .Q(\REGS[26][27] ) );
  DLH_X1 \REGS_reg[26][26]  ( .G(n372), .D(n18), .Q(\REGS[26][26] ) );
  DLH_X1 \REGS_reg[26][25]  ( .G(n372), .D(n21), .Q(\REGS[26][25] ) );
  DLH_X1 \REGS_reg[26][24]  ( .G(n372), .D(n24), .Q(\REGS[26][24] ) );
  DLH_X1 \REGS_reg[26][23]  ( .G(n372), .D(n27), .Q(\REGS[26][23] ) );
  DLH_X1 \REGS_reg[26][22]  ( .G(n372), .D(n30), .Q(\REGS[26][22] ) );
  DLH_X1 \REGS_reg[26][21]  ( .G(n371), .D(n33), .Q(\REGS[26][21] ) );
  DLH_X1 \REGS_reg[26][20]  ( .G(n371), .D(n36), .Q(\REGS[26][20] ) );
  DLH_X1 \REGS_reg[26][19]  ( .G(n371), .D(n39), .Q(\REGS[26][19] ) );
  DLH_X1 \REGS_reg[26][18]  ( .G(n371), .D(n42), .Q(\REGS[26][18] ) );
  DLH_X1 \REGS_reg[26][17]  ( .G(n371), .D(n45), .Q(\REGS[26][17] ) );
  DLH_X1 \REGS_reg[26][16]  ( .G(n371), .D(n48), .Q(\REGS[26][16] ) );
  DLH_X1 \REGS_reg[26][15]  ( .G(n371), .D(n51), .Q(\REGS[26][15] ) );
  DLH_X1 \REGS_reg[26][14]  ( .G(n371), .D(n54), .Q(\REGS[26][14] ) );
  DLH_X1 \REGS_reg[26][13]  ( .G(n371), .D(n57), .Q(\REGS[26][13] ) );
  DLH_X1 \REGS_reg[26][12]  ( .G(n371), .D(n60), .Q(\REGS[26][12] ) );
  DLH_X1 \REGS_reg[26][11]  ( .G(n371), .D(n63), .Q(\REGS[26][11] ) );
  DLH_X1 \REGS_reg[26][10]  ( .G(n370), .D(n66), .Q(\REGS[26][10] ) );
  DLH_X1 \REGS_reg[26][9]  ( .G(n370), .D(n69), .Q(\REGS[26][9] ) );
  DLH_X1 \REGS_reg[26][8]  ( .G(n370), .D(n72), .Q(\REGS[26][8] ) );
  DLH_X1 \REGS_reg[26][7]  ( .G(n370), .D(n75), .Q(\REGS[26][7] ) );
  DLH_X1 \REGS_reg[26][6]  ( .G(n370), .D(n78), .Q(\REGS[26][6] ) );
  DLH_X1 \REGS_reg[26][5]  ( .G(n370), .D(n81), .Q(\REGS[26][5] ) );
  DLH_X1 \REGS_reg[26][4]  ( .G(n370), .D(n84), .Q(\REGS[26][4] ) );
  DLH_X1 \REGS_reg[26][3]  ( .G(n370), .D(n87), .Q(\REGS[26][3] ) );
  DLH_X1 \REGS_reg[26][2]  ( .G(n370), .D(n90), .Q(\REGS[26][2] ) );
  DLH_X1 \REGS_reg[26][1]  ( .G(n370), .D(n93), .Q(\REGS[26][1] ) );
  DLH_X1 \REGS_reg[26][0]  ( .G(n370), .D(n96), .Q(\REGS[26][0] ) );
  DLH_X1 \REGS_reg[27][31]  ( .G(n375), .D(n3), .Q(\REGS[27][31] ) );
  DLH_X1 \REGS_reg[27][30]  ( .G(n375), .D(n6), .Q(\REGS[27][30] ) );
  DLH_X1 \REGS_reg[27][29]  ( .G(n375), .D(n9), .Q(\REGS[27][29] ) );
  DLH_X1 \REGS_reg[27][28]  ( .G(n375), .D(n12), .Q(\REGS[27][28] ) );
  DLH_X1 \REGS_reg[27][27]  ( .G(n375), .D(n15), .Q(\REGS[27][27] ) );
  DLH_X1 \REGS_reg[27][26]  ( .G(n375), .D(n18), .Q(\REGS[27][26] ) );
  DLH_X1 \REGS_reg[27][25]  ( .G(n375), .D(n21), .Q(\REGS[27][25] ) );
  DLH_X1 \REGS_reg[27][24]  ( .G(n375), .D(n24), .Q(\REGS[27][24] ) );
  DLH_X1 \REGS_reg[27][23]  ( .G(n375), .D(n27), .Q(\REGS[27][23] ) );
  DLH_X1 \REGS_reg[27][22]  ( .G(n375), .D(n30), .Q(\REGS[27][22] ) );
  DLH_X1 \REGS_reg[27][21]  ( .G(n374), .D(n33), .Q(\REGS[27][21] ) );
  DLH_X1 \REGS_reg[27][20]  ( .G(n374), .D(n36), .Q(\REGS[27][20] ) );
  DLH_X1 \REGS_reg[27][19]  ( .G(n374), .D(n39), .Q(\REGS[27][19] ) );
  DLH_X1 \REGS_reg[27][18]  ( .G(n374), .D(n42), .Q(\REGS[27][18] ) );
  DLH_X1 \REGS_reg[27][17]  ( .G(n374), .D(n45), .Q(\REGS[27][17] ) );
  DLH_X1 \REGS_reg[27][16]  ( .G(n374), .D(n48), .Q(\REGS[27][16] ) );
  DLH_X1 \REGS_reg[27][15]  ( .G(n374), .D(n51), .Q(\REGS[27][15] ) );
  DLH_X1 \REGS_reg[27][14]  ( .G(n374), .D(n54), .Q(\REGS[27][14] ) );
  DLH_X1 \REGS_reg[27][13]  ( .G(n374), .D(n57), .Q(\REGS[27][13] ) );
  DLH_X1 \REGS_reg[27][12]  ( .G(n374), .D(n60), .Q(\REGS[27][12] ) );
  DLH_X1 \REGS_reg[27][11]  ( .G(n374), .D(n63), .Q(\REGS[27][11] ) );
  DLH_X1 \REGS_reg[27][10]  ( .G(n373), .D(n66), .Q(\REGS[27][10] ) );
  DLH_X1 \REGS_reg[27][9]  ( .G(n373), .D(n69), .Q(\REGS[27][9] ) );
  DLH_X1 \REGS_reg[27][8]  ( .G(n373), .D(n72), .Q(\REGS[27][8] ) );
  DLH_X1 \REGS_reg[27][7]  ( .G(n373), .D(n75), .Q(\REGS[27][7] ) );
  DLH_X1 \REGS_reg[27][6]  ( .G(n373), .D(n78), .Q(\REGS[27][6] ) );
  DLH_X1 \REGS_reg[27][5]  ( .G(n373), .D(n81), .Q(\REGS[27][5] ) );
  DLH_X1 \REGS_reg[27][4]  ( .G(n373), .D(n84), .Q(\REGS[27][4] ) );
  DLH_X1 \REGS_reg[27][3]  ( .G(n373), .D(n87), .Q(\REGS[27][3] ) );
  DLH_X1 \REGS_reg[27][2]  ( .G(n373), .D(n90), .Q(\REGS[27][2] ) );
  DLH_X1 \REGS_reg[27][1]  ( .G(n373), .D(n93), .Q(\REGS[27][1] ) );
  DLH_X1 \REGS_reg[27][0]  ( .G(n373), .D(n96), .Q(\REGS[27][0] ) );
  DLH_X1 \REGS_reg[28][31]  ( .G(n378), .D(n3), .Q(\REGS[28][31] ) );
  DLH_X1 \REGS_reg[28][30]  ( .G(n378), .D(n6), .Q(\REGS[28][30] ) );
  DLH_X1 \REGS_reg[28][29]  ( .G(n378), .D(n9), .Q(\REGS[28][29] ) );
  DLH_X1 \REGS_reg[28][28]  ( .G(n378), .D(n12), .Q(\REGS[28][28] ) );
  DLH_X1 \REGS_reg[28][27]  ( .G(n378), .D(n15), .Q(\REGS[28][27] ) );
  DLH_X1 \REGS_reg[28][26]  ( .G(n378), .D(n18), .Q(\REGS[28][26] ) );
  DLH_X1 \REGS_reg[28][25]  ( .G(n378), .D(n21), .Q(\REGS[28][25] ) );
  DLH_X1 \REGS_reg[28][24]  ( .G(n378), .D(n24), .Q(\REGS[28][24] ) );
  DLH_X1 \REGS_reg[28][23]  ( .G(n378), .D(n27), .Q(\REGS[28][23] ) );
  DLH_X1 \REGS_reg[28][22]  ( .G(n378), .D(n30), .Q(\REGS[28][22] ) );
  DLH_X1 \REGS_reg[28][21]  ( .G(n377), .D(n33), .Q(\REGS[28][21] ) );
  DLH_X1 \REGS_reg[28][20]  ( .G(n377), .D(n36), .Q(\REGS[28][20] ) );
  DLH_X1 \REGS_reg[28][19]  ( .G(n377), .D(n39), .Q(\REGS[28][19] ) );
  DLH_X1 \REGS_reg[28][18]  ( .G(n377), .D(n42), .Q(\REGS[28][18] ) );
  DLH_X1 \REGS_reg[28][17]  ( .G(n377), .D(n45), .Q(\REGS[28][17] ) );
  DLH_X1 \REGS_reg[28][16]  ( .G(n377), .D(n48), .Q(\REGS[28][16] ) );
  DLH_X1 \REGS_reg[28][15]  ( .G(n377), .D(n51), .Q(\REGS[28][15] ) );
  DLH_X1 \REGS_reg[28][14]  ( .G(n377), .D(n54), .Q(\REGS[28][14] ) );
  DLH_X1 \REGS_reg[28][13]  ( .G(n377), .D(n57), .Q(\REGS[28][13] ) );
  DLH_X1 \REGS_reg[28][12]  ( .G(n377), .D(n60), .Q(\REGS[28][12] ) );
  DLH_X1 \REGS_reg[28][11]  ( .G(n377), .D(n63), .Q(\REGS[28][11] ) );
  DLH_X1 \REGS_reg[28][10]  ( .G(n376), .D(n66), .Q(\REGS[28][10] ) );
  DLH_X1 \REGS_reg[28][9]  ( .G(n376), .D(n69), .Q(\REGS[28][9] ) );
  DLH_X1 \REGS_reg[28][8]  ( .G(n376), .D(n72), .Q(\REGS[28][8] ) );
  DLH_X1 \REGS_reg[28][7]  ( .G(n376), .D(n75), .Q(\REGS[28][7] ) );
  DLH_X1 \REGS_reg[28][6]  ( .G(n376), .D(n78), .Q(\REGS[28][6] ) );
  DLH_X1 \REGS_reg[28][5]  ( .G(n376), .D(n81), .Q(\REGS[28][5] ) );
  DLH_X1 \REGS_reg[28][4]  ( .G(n376), .D(n84), .Q(\REGS[28][4] ) );
  DLH_X1 \REGS_reg[28][3]  ( .G(n376), .D(n87), .Q(\REGS[28][3] ) );
  DLH_X1 \REGS_reg[28][2]  ( .G(n376), .D(n90), .Q(\REGS[28][2] ) );
  DLH_X1 \REGS_reg[28][1]  ( .G(n376), .D(n93), .Q(\REGS[28][1] ) );
  DLH_X1 \REGS_reg[28][0]  ( .G(n376), .D(n96), .Q(\REGS[28][0] ) );
  DLH_X1 \REGS_reg[29][31]  ( .G(n381), .D(n3), .Q(\REGS[29][31] ) );
  DLH_X1 \REGS_reg[29][30]  ( .G(n381), .D(n6), .Q(\REGS[29][30] ) );
  DLH_X1 \REGS_reg[29][29]  ( .G(n381), .D(n9), .Q(\REGS[29][29] ) );
  DLH_X1 \REGS_reg[29][28]  ( .G(n381), .D(n12), .Q(\REGS[29][28] ) );
  DLH_X1 \REGS_reg[29][27]  ( .G(n381), .D(n15), .Q(\REGS[29][27] ) );
  DLH_X1 \REGS_reg[29][26]  ( .G(n381), .D(n18), .Q(\REGS[29][26] ) );
  DLH_X1 \REGS_reg[29][25]  ( .G(n381), .D(n21), .Q(\REGS[29][25] ) );
  DLH_X1 \REGS_reg[29][24]  ( .G(n381), .D(n24), .Q(\REGS[29][24] ) );
  DLH_X1 \REGS_reg[29][23]  ( .G(n381), .D(n27), .Q(\REGS[29][23] ) );
  DLH_X1 \REGS_reg[29][22]  ( .G(n381), .D(n30), .Q(\REGS[29][22] ) );
  DLH_X1 \REGS_reg[29][21]  ( .G(n380), .D(n33), .Q(\REGS[29][21] ) );
  DLH_X1 \REGS_reg[29][20]  ( .G(n380), .D(n36), .Q(\REGS[29][20] ) );
  DLH_X1 \REGS_reg[29][19]  ( .G(n380), .D(n39), .Q(\REGS[29][19] ) );
  DLH_X1 \REGS_reg[29][18]  ( .G(n380), .D(n42), .Q(\REGS[29][18] ) );
  DLH_X1 \REGS_reg[29][17]  ( .G(n380), .D(n45), .Q(\REGS[29][17] ) );
  DLH_X1 \REGS_reg[29][16]  ( .G(n380), .D(n48), .Q(\REGS[29][16] ) );
  DLH_X1 \REGS_reg[29][15]  ( .G(n380), .D(n51), .Q(\REGS[29][15] ) );
  DLH_X1 \REGS_reg[29][14]  ( .G(n380), .D(n54), .Q(\REGS[29][14] ) );
  DLH_X1 \REGS_reg[29][13]  ( .G(n380), .D(n57), .Q(\REGS[29][13] ) );
  DLH_X1 \REGS_reg[29][12]  ( .G(n380), .D(n60), .Q(\REGS[29][12] ) );
  DLH_X1 \REGS_reg[29][11]  ( .G(n380), .D(n63), .Q(\REGS[29][11] ) );
  DLH_X1 \REGS_reg[29][10]  ( .G(n379), .D(n66), .Q(\REGS[29][10] ) );
  DLH_X1 \REGS_reg[29][9]  ( .G(n379), .D(n69), .Q(\REGS[29][9] ) );
  DLH_X1 \REGS_reg[29][8]  ( .G(n379), .D(n72), .Q(\REGS[29][8] ) );
  DLH_X1 \REGS_reg[29][7]  ( .G(n379), .D(n75), .Q(\REGS[29][7] ) );
  DLH_X1 \REGS_reg[29][6]  ( .G(n379), .D(n78), .Q(\REGS[29][6] ) );
  DLH_X1 \REGS_reg[29][5]  ( .G(n379), .D(n81), .Q(\REGS[29][5] ) );
  DLH_X1 \REGS_reg[29][4]  ( .G(n379), .D(n84), .Q(\REGS[29][4] ) );
  DLH_X1 \REGS_reg[29][3]  ( .G(n379), .D(n87), .Q(\REGS[29][3] ) );
  DLH_X1 \REGS_reg[29][2]  ( .G(n379), .D(n90), .Q(\REGS[29][2] ) );
  DLH_X1 \REGS_reg[29][1]  ( .G(n379), .D(n93), .Q(\REGS[29][1] ) );
  DLH_X1 \REGS_reg[29][0]  ( .G(n379), .D(n96), .Q(\REGS[29][0] ) );
  DLH_X1 \REGS_reg[30][31]  ( .G(n384), .D(n3), .Q(\REGS[30][31] ) );
  DLH_X1 \REGS_reg[30][30]  ( .G(n384), .D(n6), .Q(\REGS[30][30] ) );
  DLH_X1 \REGS_reg[30][29]  ( .G(n384), .D(n9), .Q(\REGS[30][29] ) );
  DLH_X1 \REGS_reg[30][28]  ( .G(n384), .D(n12), .Q(\REGS[30][28] ) );
  DLH_X1 \REGS_reg[30][27]  ( .G(n384), .D(n15), .Q(\REGS[30][27] ) );
  DLH_X1 \REGS_reg[30][26]  ( .G(n384), .D(n18), .Q(\REGS[30][26] ) );
  DLH_X1 \REGS_reg[30][25]  ( .G(n384), .D(n21), .Q(\REGS[30][25] ) );
  DLH_X1 \REGS_reg[30][24]  ( .G(n384), .D(n24), .Q(\REGS[30][24] ) );
  DLH_X1 \REGS_reg[30][23]  ( .G(n384), .D(n27), .Q(\REGS[30][23] ) );
  DLH_X1 \REGS_reg[30][22]  ( .G(n384), .D(n30), .Q(\REGS[30][22] ) );
  DLH_X1 \REGS_reg[30][21]  ( .G(n383), .D(n33), .Q(\REGS[30][21] ) );
  DLH_X1 \REGS_reg[30][20]  ( .G(n383), .D(n36), .Q(\REGS[30][20] ) );
  DLH_X1 \REGS_reg[30][19]  ( .G(n383), .D(n39), .Q(\REGS[30][19] ) );
  DLH_X1 \REGS_reg[30][18]  ( .G(n383), .D(n42), .Q(\REGS[30][18] ) );
  DLH_X1 \REGS_reg[30][17]  ( .G(n383), .D(n45), .Q(\REGS[30][17] ) );
  DLH_X1 \REGS_reg[30][16]  ( .G(n383), .D(n48), .Q(\REGS[30][16] ) );
  DLH_X1 \REGS_reg[30][15]  ( .G(n383), .D(n51), .Q(\REGS[30][15] ) );
  DLH_X1 \REGS_reg[30][14]  ( .G(n383), .D(n54), .Q(\REGS[30][14] ) );
  DLH_X1 \REGS_reg[30][13]  ( .G(n383), .D(n57), .Q(\REGS[30][13] ) );
  DLH_X1 \REGS_reg[30][12]  ( .G(n383), .D(n60), .Q(\REGS[30][12] ) );
  DLH_X1 \REGS_reg[30][11]  ( .G(n383), .D(n63), .Q(\REGS[30][11] ) );
  DLH_X1 \REGS_reg[30][10]  ( .G(n382), .D(n66), .Q(\REGS[30][10] ) );
  DLH_X1 \REGS_reg[30][9]  ( .G(n382), .D(n69), .Q(\REGS[30][9] ) );
  DLH_X1 \REGS_reg[30][8]  ( .G(n382), .D(n72), .Q(\REGS[30][8] ) );
  DLH_X1 \REGS_reg[30][7]  ( .G(n382), .D(n75), .Q(\REGS[30][7] ) );
  DLH_X1 \REGS_reg[30][6]  ( .G(n382), .D(n78), .Q(\REGS[30][6] ) );
  DLH_X1 \REGS_reg[30][5]  ( .G(n382), .D(n81), .Q(\REGS[30][5] ) );
  DLH_X1 \REGS_reg[30][4]  ( .G(n382), .D(n84), .Q(\REGS[30][4] ) );
  DLH_X1 \REGS_reg[30][3]  ( .G(n382), .D(n87), .Q(\REGS[30][3] ) );
  DLH_X1 \REGS_reg[30][2]  ( .G(n382), .D(n90), .Q(\REGS[30][2] ) );
  DLH_X1 \REGS_reg[30][1]  ( .G(n382), .D(n93), .Q(\REGS[30][1] ) );
  DLH_X1 \REGS_reg[30][0]  ( .G(n382), .D(n96), .Q(\REGS[30][0] ) );
  DLH_X1 \REGS_reg[31][31]  ( .G(n387), .D(n3), .Q(\REGS[31][31] ) );
  DLL_X1 \DATA_OUT1_reg[31]  ( .D(N79), .GN(n392), .Q(DATA_OUT1[31]) );
  DLL_X1 \DATA_OUT2_reg[31]  ( .D(N176), .GN(n392), .Q(DATA_OUT2[31]) );
  DLH_X1 \REGS_reg[31][30]  ( .G(n387), .D(n6), .Q(\REGS[31][30] ) );
  DLL_X1 \DATA_OUT1_reg[30]  ( .D(N80), .GN(n392), .Q(DATA_OUT1[30]) );
  DLL_X1 \DATA_OUT2_reg[30]  ( .D(N177), .GN(n392), .Q(DATA_OUT2[30]) );
  DLH_X1 \REGS_reg[31][29]  ( .G(n387), .D(n9), .Q(\REGS[31][29] ) );
  DLL_X1 \DATA_OUT1_reg[29]  ( .D(N81), .GN(n392), .Q(DATA_OUT1[29]) );
  DLL_X1 \DATA_OUT2_reg[29]  ( .D(N178), .GN(n392), .Q(DATA_OUT2[29]) );
  DLH_X1 \REGS_reg[31][28]  ( .G(n387), .D(n12), .Q(\REGS[31][28] ) );
  DLL_X1 \DATA_OUT1_reg[28]  ( .D(N82), .GN(n392), .Q(DATA_OUT1[28]) );
  DLL_X1 \DATA_OUT2_reg[28]  ( .D(N179), .GN(n392), .Q(DATA_OUT2[28]) );
  DLH_X1 \REGS_reg[31][27]  ( .G(n387), .D(n15), .Q(\REGS[31][27] ) );
  DLL_X1 \DATA_OUT1_reg[27]  ( .D(N83), .GN(n392), .Q(DATA_OUT1[27]) );
  DLL_X1 \DATA_OUT2_reg[27]  ( .D(N180), .GN(n392), .Q(DATA_OUT2[27]) );
  DLH_X1 \REGS_reg[31][26]  ( .G(n387), .D(n18), .Q(\REGS[31][26] ) );
  DLL_X1 \DATA_OUT1_reg[26]  ( .D(N84), .GN(n392), .Q(DATA_OUT1[26]) );
  DLL_X1 \DATA_OUT2_reg[26]  ( .D(N181), .GN(n392), .Q(DATA_OUT2[26]) );
  DLH_X1 \REGS_reg[31][25]  ( .G(n387), .D(n21), .Q(\REGS[31][25] ) );
  DLL_X1 \DATA_OUT1_reg[25]  ( .D(N85), .GN(n393), .Q(DATA_OUT1[25]) );
  DLL_X1 \DATA_OUT2_reg[25]  ( .D(N182), .GN(n393), .Q(DATA_OUT2[25]) );
  DLH_X1 \REGS_reg[31][24]  ( .G(n387), .D(n24), .Q(\REGS[31][24] ) );
  DLL_X1 \DATA_OUT1_reg[24]  ( .D(N86), .GN(n393), .Q(DATA_OUT1[24]) );
  DLL_X1 \DATA_OUT2_reg[24]  ( .D(N183), .GN(n394), .Q(DATA_OUT2[24]) );
  DLH_X1 \REGS_reg[31][23]  ( .G(n387), .D(n27), .Q(\REGS[31][23] ) );
  DLL_X1 \DATA_OUT1_reg[23]  ( .D(N87), .GN(n393), .Q(DATA_OUT1[23]) );
  DLL_X1 \DATA_OUT2_reg[23]  ( .D(N184), .GN(n393), .Q(DATA_OUT2[23]) );
  DLH_X1 \REGS_reg[31][22]  ( .G(n387), .D(n30), .Q(\REGS[31][22] ) );
  DLL_X1 \DATA_OUT1_reg[22]  ( .D(N88), .GN(n393), .Q(DATA_OUT1[22]) );
  DLL_X1 \DATA_OUT2_reg[22]  ( .D(N185), .GN(n393), .Q(DATA_OUT2[22]) );
  DLH_X1 \REGS_reg[31][21]  ( .G(n386), .D(n33), .Q(\REGS[31][21] ) );
  DLL_X1 \DATA_OUT1_reg[21]  ( .D(N89), .GN(n393), .Q(DATA_OUT1[21]) );
  DLL_X1 \DATA_OUT2_reg[21]  ( .D(N186), .GN(n393), .Q(DATA_OUT2[21]) );
  DLH_X1 \REGS_reg[31][20]  ( .G(n386), .D(n36), .Q(\REGS[31][20] ) );
  DLL_X1 \DATA_OUT1_reg[20]  ( .D(N90), .GN(n393), .Q(DATA_OUT1[20]) );
  DLL_X1 \DATA_OUT2_reg[20]  ( .D(N187), .GN(n393), .Q(DATA_OUT2[20]) );
  DLH_X1 \REGS_reg[31][19]  ( .G(n386), .D(n39), .Q(\REGS[31][19] ) );
  DLL_X1 \DATA_OUT1_reg[19]  ( .D(N91), .GN(n393), .Q(DATA_OUT1[19]) );
  DLL_X1 \DATA_OUT2_reg[19]  ( .D(N188), .GN(n394), .Q(DATA_OUT2[19]) );
  DLH_X1 \REGS_reg[31][18]  ( .G(n386), .D(n42), .Q(\REGS[31][18] ) );
  DLL_X1 \DATA_OUT1_reg[18]  ( .D(N92), .GN(n394), .Q(DATA_OUT1[18]) );
  DLL_X1 \DATA_OUT2_reg[18]  ( .D(N189), .GN(n394), .Q(DATA_OUT2[18]) );
  DLH_X1 \REGS_reg[31][17]  ( .G(n386), .D(n45), .Q(\REGS[31][17] ) );
  DLL_X1 \DATA_OUT1_reg[17]  ( .D(N93), .GN(n394), .Q(DATA_OUT1[17]) );
  DLL_X1 \DATA_OUT2_reg[17]  ( .D(N190), .GN(n394), .Q(DATA_OUT2[17]) );
  DLH_X1 \REGS_reg[31][16]  ( .G(n386), .D(n48), .Q(\REGS[31][16] ) );
  DLL_X1 \DATA_OUT1_reg[16]  ( .D(N94), .GN(n394), .Q(DATA_OUT1[16]) );
  DLL_X1 \DATA_OUT2_reg[16]  ( .D(N191), .GN(n394), .Q(DATA_OUT2[16]) );
  DLH_X1 \REGS_reg[31][15]  ( .G(n386), .D(n51), .Q(\REGS[31][15] ) );
  DLL_X1 \DATA_OUT1_reg[15]  ( .D(N95), .GN(n394), .Q(DATA_OUT1[15]) );
  DLL_X1 \DATA_OUT2_reg[15]  ( .D(N192), .GN(n394), .Q(DATA_OUT2[15]) );
  DLH_X1 \REGS_reg[31][14]  ( .G(n386), .D(n54), .Q(\REGS[31][14] ) );
  DLL_X1 \DATA_OUT1_reg[14]  ( .D(N96), .GN(n394), .Q(DATA_OUT1[14]) );
  DLL_X1 \DATA_OUT2_reg[14]  ( .D(N193), .GN(n394), .Q(DATA_OUT2[14]) );
  DLH_X1 \REGS_reg[31][13]  ( .G(n386), .D(n57), .Q(\REGS[31][13] ) );
  DLL_X1 \DATA_OUT1_reg[13]  ( .D(N97), .GN(n395), .Q(DATA_OUT1[13]) );
  DLL_X1 \DATA_OUT2_reg[13]  ( .D(N194), .GN(n395), .Q(DATA_OUT2[13]) );
  DLH_X1 \REGS_reg[31][12]  ( .G(n386), .D(n60), .Q(\REGS[31][12] ) );
  DLL_X1 \DATA_OUT1_reg[12]  ( .D(N98), .GN(n395), .Q(DATA_OUT1[12]) );
  DLL_X1 \DATA_OUT2_reg[12]  ( .D(N195), .GN(n395), .Q(DATA_OUT2[12]) );
  DLH_X1 \REGS_reg[31][11]  ( .G(n386), .D(n63), .Q(\REGS[31][11] ) );
  DLL_X1 \DATA_OUT1_reg[11]  ( .D(N99), .GN(n395), .Q(DATA_OUT1[11]) );
  DLL_X1 \DATA_OUT2_reg[11]  ( .D(N196), .GN(n395), .Q(DATA_OUT2[11]) );
  DLH_X1 \REGS_reg[31][10]  ( .G(n385), .D(n66), .Q(\REGS[31][10] ) );
  DLL_X1 \DATA_OUT2_reg[10]  ( .D(N197), .GN(n395), .Q(DATA_OUT2[10]) );
  DLL_X1 \DATA_OUT1_reg[10]  ( .D(N100), .GN(n395), .Q(DATA_OUT1[10]) );
  DLH_X1 \REGS_reg[31][9]  ( .G(n385), .D(n69), .Q(\REGS[31][9] ) );
  DLL_X1 \DATA_OUT2_reg[9]  ( .D(N198), .GN(n395), .Q(DATA_OUT2[9]) );
  DLL_X1 \DATA_OUT1_reg[9]  ( .D(N101), .GN(n395), .Q(DATA_OUT1[9]) );
  DLH_X1 \REGS_reg[31][8]  ( .G(n385), .D(n72), .Q(\REGS[31][8] ) );
  DLL_X1 \DATA_OUT2_reg[8]  ( .D(N199), .GN(n395), .Q(DATA_OUT2[8]) );
  DLL_X1 \DATA_OUT1_reg[8]  ( .D(N102), .GN(n395), .Q(DATA_OUT1[8]) );
  DLH_X1 \REGS_reg[31][7]  ( .G(n385), .D(n75), .Q(\REGS[31][7] ) );
  DLL_X1 \DATA_OUT2_reg[7]  ( .D(N200), .GN(n396), .Q(DATA_OUT2[7]) );
  DLL_X1 \DATA_OUT1_reg[7]  ( .D(N103), .GN(n396), .Q(DATA_OUT1[7]) );
  DLH_X1 \REGS_reg[31][6]  ( .G(n385), .D(n78), .Q(\REGS[31][6] ) );
  DLL_X1 \DATA_OUT2_reg[6]  ( .D(N201), .GN(n396), .Q(DATA_OUT2[6]) );
  DLL_X1 \DATA_OUT1_reg[6]  ( .D(N104), .GN(n396), .Q(DATA_OUT1[6]) );
  DLH_X1 \REGS_reg[31][5]  ( .G(n385), .D(n81), .Q(\REGS[31][5] ) );
  DLL_X1 \DATA_OUT2_reg[5]  ( .D(N202), .GN(n396), .Q(DATA_OUT2[5]) );
  DLL_X1 \DATA_OUT1_reg[5]  ( .D(N105), .GN(n396), .Q(DATA_OUT1[5]) );
  DLH_X1 \REGS_reg[31][4]  ( .G(n385), .D(n84), .Q(\REGS[31][4] ) );
  DLL_X1 \DATA_OUT2_reg[4]  ( .D(N203), .GN(n396), .Q(DATA_OUT2[4]) );
  DLL_X1 \DATA_OUT1_reg[4]  ( .D(N106), .GN(n396), .Q(DATA_OUT1[4]) );
  DLH_X1 \REGS_reg[31][3]  ( .G(n385), .D(n87), .Q(\REGS[31][3] ) );
  DLL_X1 \DATA_OUT2_reg[3]  ( .D(N204), .GN(n396), .Q(DATA_OUT2[3]) );
  DLL_X1 \DATA_OUT1_reg[3]  ( .D(N107), .GN(n396), .Q(DATA_OUT1[3]) );
  DLH_X1 \REGS_reg[31][2]  ( .G(n385), .D(n90), .Q(\REGS[31][2] ) );
  DLL_X1 \DATA_OUT2_reg[2]  ( .D(N205), .GN(n396), .Q(DATA_OUT2[2]) );
  DLL_X1 \DATA_OUT1_reg[2]  ( .D(N108), .GN(n396), .Q(DATA_OUT1[2]) );
  DLH_X1 \REGS_reg[31][1]  ( .G(n385), .D(n93), .Q(\REGS[31][1] ) );
  DLL_X1 \DATA_OUT2_reg[1]  ( .D(N206), .GN(n397), .Q(DATA_OUT2[1]) );
  DLL_X1 \DATA_OUT1_reg[1]  ( .D(N109), .GN(n397), .Q(DATA_OUT1[1]) );
  DLH_X1 \REGS_reg[31][0]  ( .G(n385), .D(n96), .Q(\REGS[31][0] ) );
  DLL_X1 \DATA_OUT2_reg[0]  ( .D(N207), .GN(n397), .Q(DATA_OUT2[0]) );
  DLL_X1 \DATA_OUT1_reg[0]  ( .D(N110), .GN(n391), .Q(DATA_OUT1[0]) );
  NAND3_X1 U1970 ( .A1(n399), .A2(n398), .A3(WE), .ZN(n1004) );
  NAND3_X1 U1971 ( .A1(WE), .A2(n398), .A3(ADDR_WR[3]), .ZN(n1012) );
  NAND3_X1 U1972 ( .A1(WE), .A2(n399), .A3(ADDR_WR[4]), .ZN(n1013) );
  NAND3_X1 U1973 ( .A1(n401), .A2(n400), .A3(n402), .ZN(n1003) );
  NAND3_X1 U1974 ( .A1(n401), .A2(n400), .A3(ADDR_WR[0]), .ZN(n1005) );
  NAND3_X1 U1975 ( .A1(n402), .A2(n400), .A3(ADDR_WR[1]), .ZN(n1006) );
  NAND3_X1 U1976 ( .A1(ADDR_WR[0]), .A2(n400), .A3(ADDR_WR[1]), .ZN(n1007) );
  NAND3_X1 U1977 ( .A1(n402), .A2(n401), .A3(ADDR_WR[2]), .ZN(n1008) );
  NAND3_X1 U1978 ( .A1(ADDR_WR[0]), .A2(n401), .A3(ADDR_WR[2]), .ZN(n1009) );
  NAND3_X1 U1979 ( .A1(ADDR_WR[1]), .A2(n402), .A3(ADDR_WR[2]), .ZN(n1010) );
  NAND3_X1 U1980 ( .A1(ADDR_WR[3]), .A2(WE), .A3(ADDR_WR[4]), .ZN(n1014) );
  NAND3_X1 U1981 ( .A1(ADDR_WR[1]), .A2(ADDR_WR[0]), .A3(ADDR_WR[2]), .ZN(
        n1011) );
  NOR2_X1 U3 ( .A1(n408), .A2(ADDR_RD2[1]), .ZN(n1618) );
  NOR2_X1 U4 ( .A1(n404), .A2(ADDR_RD1[1]), .ZN(n1832) );
  NOR2_X1 U5 ( .A1(ADDR_RD2[1]), .A2(ADDR_RD2[2]), .ZN(n1615) );
  NOR2_X1 U6 ( .A1(ADDR_RD1[1]), .A2(ADDR_RD1[2]), .ZN(n1829) );
  BUF_X1 U7 ( .A(n574), .Z(n272) );
  BUF_X1 U8 ( .A(n598), .Z(n224) );
  BUF_X1 U9 ( .A(n608), .Z(n200) );
  BUF_X1 U10 ( .A(n574), .Z(n271) );
  BUF_X1 U11 ( .A(n598), .Z(n223) );
  BUF_X1 U12 ( .A(n608), .Z(n199) );
  BUF_X1 U13 ( .A(n1030), .Z(n169) );
  BUF_X1 U14 ( .A(n1054), .Z(n121) );
  BUF_X1 U15 ( .A(n1064), .Z(n97) );
  BUF_X1 U16 ( .A(n1030), .Z(n170) );
  BUF_X1 U17 ( .A(n1054), .Z(n122) );
  BUF_X1 U18 ( .A(n1064), .Z(n98) );
  BUF_X1 U19 ( .A(n1037), .Z(n151) );
  BUF_X1 U20 ( .A(n1037), .Z(n152) );
  BUF_X1 U21 ( .A(n574), .Z(n273) );
  BUF_X1 U22 ( .A(n598), .Z(n225) );
  BUF_X1 U23 ( .A(n608), .Z(n201) );
  BUF_X1 U24 ( .A(n581), .Z(n254) );
  BUF_X1 U25 ( .A(n581), .Z(n253) );
  BUF_X1 U26 ( .A(n1037), .Z(n153) );
  BUF_X1 U27 ( .A(n581), .Z(n255) );
  BUF_X1 U28 ( .A(n1030), .Z(n171) );
  BUF_X1 U29 ( .A(n1054), .Z(n123) );
  BUF_X1 U30 ( .A(n1064), .Z(n99) );
  INV_X1 U31 ( .A(n391), .ZN(n390) );
  INV_X1 U32 ( .A(n391), .ZN(n388) );
  INV_X1 U33 ( .A(n391), .ZN(n389) );
  BUF_X1 U34 ( .A(n1024), .Z(n185) );
  BUF_X1 U35 ( .A(n1029), .Z(n173) );
  BUF_X1 U36 ( .A(n1034), .Z(n161) );
  BUF_X1 U37 ( .A(n1039), .Z(n149) );
  BUF_X1 U38 ( .A(n1048), .Z(n137) );
  BUF_X1 U39 ( .A(n1053), .Z(n125) );
  BUF_X1 U40 ( .A(n1058), .Z(n113) );
  BUF_X1 U41 ( .A(n1063), .Z(n101) );
  BUF_X1 U42 ( .A(n568), .Z(n287) );
  BUF_X1 U43 ( .A(n573), .Z(n275) );
  BUF_X1 U44 ( .A(n578), .Z(n263) );
  BUF_X1 U45 ( .A(n583), .Z(n251) );
  BUF_X1 U46 ( .A(n592), .Z(n239) );
  BUF_X1 U47 ( .A(n597), .Z(n227) );
  BUF_X1 U48 ( .A(n602), .Z(n215) );
  BUF_X1 U49 ( .A(n607), .Z(n203) );
  BUF_X1 U50 ( .A(n568), .Z(n286) );
  BUF_X1 U51 ( .A(n573), .Z(n274) );
  BUF_X1 U52 ( .A(n578), .Z(n262) );
  BUF_X1 U53 ( .A(n583), .Z(n250) );
  BUF_X1 U54 ( .A(n592), .Z(n238) );
  BUF_X1 U55 ( .A(n597), .Z(n226) );
  BUF_X1 U56 ( .A(n602), .Z(n214) );
  BUF_X1 U57 ( .A(n607), .Z(n202) );
  BUF_X1 U58 ( .A(n565), .Z(n293) );
  BUF_X1 U59 ( .A(n570), .Z(n281) );
  BUF_X1 U60 ( .A(n575), .Z(n269) );
  BUF_X1 U61 ( .A(n580), .Z(n257) );
  BUF_X1 U62 ( .A(n589), .Z(n245) );
  BUF_X1 U63 ( .A(n594), .Z(n233) );
  BUF_X1 U64 ( .A(n599), .Z(n221) );
  BUF_X1 U65 ( .A(n604), .Z(n209) );
  BUF_X1 U66 ( .A(n565), .Z(n292) );
  BUF_X1 U67 ( .A(n570), .Z(n280) );
  BUF_X1 U68 ( .A(n575), .Z(n268) );
  BUF_X1 U69 ( .A(n580), .Z(n256) );
  BUF_X1 U70 ( .A(n589), .Z(n244) );
  BUF_X1 U71 ( .A(n594), .Z(n232) );
  BUF_X1 U72 ( .A(n599), .Z(n220) );
  BUF_X1 U73 ( .A(n604), .Z(n208) );
  BUF_X1 U74 ( .A(n1021), .Z(n191) );
  BUF_X1 U75 ( .A(n1045), .Z(n143) );
  BUF_X1 U76 ( .A(n1055), .Z(n119) );
  BUF_X1 U77 ( .A(n1026), .Z(n179) );
  BUF_X1 U78 ( .A(n1050), .Z(n131) );
  BUF_X1 U79 ( .A(n1060), .Z(n107) );
  BUF_X1 U80 ( .A(n1031), .Z(n167) );
  BUF_X1 U81 ( .A(n1036), .Z(n155) );
  BUF_X1 U82 ( .A(n1024), .Z(n184) );
  BUF_X1 U83 ( .A(n1029), .Z(n172) );
  BUF_X1 U84 ( .A(n1034), .Z(n160) );
  BUF_X1 U85 ( .A(n1039), .Z(n148) );
  BUF_X1 U86 ( .A(n1048), .Z(n136) );
  BUF_X1 U87 ( .A(n1053), .Z(n124) );
  BUF_X1 U88 ( .A(n1058), .Z(n112) );
  BUF_X1 U89 ( .A(n1063), .Z(n100) );
  BUF_X1 U90 ( .A(n1021), .Z(n190) );
  BUF_X1 U91 ( .A(n1045), .Z(n142) );
  BUF_X1 U92 ( .A(n1055), .Z(n118) );
  BUF_X1 U93 ( .A(n1026), .Z(n178) );
  BUF_X1 U94 ( .A(n1050), .Z(n130) );
  BUF_X1 U95 ( .A(n1060), .Z(n106) );
  BUF_X1 U96 ( .A(n1031), .Z(n166) );
  BUF_X1 U97 ( .A(n1036), .Z(n154) );
  BUF_X1 U98 ( .A(n569), .Z(n284) );
  BUF_X1 U99 ( .A(n579), .Z(n260) );
  BUF_X1 U100 ( .A(n584), .Z(n248) );
  BUF_X1 U101 ( .A(n593), .Z(n236) );
  BUF_X1 U102 ( .A(n603), .Z(n212) );
  BUF_X1 U103 ( .A(n569), .Z(n283) );
  BUF_X1 U104 ( .A(n579), .Z(n259) );
  BUF_X1 U105 ( .A(n584), .Z(n247) );
  BUF_X1 U106 ( .A(n593), .Z(n235) );
  BUF_X1 U107 ( .A(n603), .Z(n211) );
  BUF_X1 U108 ( .A(n969), .Z(n198) );
  BUF_X1 U109 ( .A(n1025), .Z(n181) );
  BUF_X1 U110 ( .A(n1035), .Z(n157) );
  BUF_X1 U111 ( .A(n1040), .Z(n145) );
  BUF_X1 U112 ( .A(n1049), .Z(n133) );
  BUF_X1 U113 ( .A(n1059), .Z(n109) );
  BUF_X1 U114 ( .A(n969), .Z(n197) );
  BUF_X1 U115 ( .A(n969), .Z(n196) );
  BUF_X1 U116 ( .A(n1025), .Z(n182) );
  BUF_X1 U117 ( .A(n1035), .Z(n158) );
  BUF_X1 U118 ( .A(n1040), .Z(n146) );
  BUF_X1 U119 ( .A(n1049), .Z(n134) );
  BUF_X1 U120 ( .A(n1059), .Z(n110) );
  BUF_X1 U121 ( .A(n1022), .Z(n187) );
  BUF_X1 U122 ( .A(n1046), .Z(n139) );
  BUF_X1 U123 ( .A(n1056), .Z(n115) );
  BUF_X1 U124 ( .A(n1027), .Z(n175) );
  BUF_X1 U125 ( .A(n1051), .Z(n127) );
  BUF_X1 U126 ( .A(n1061), .Z(n103) );
  BUF_X1 U127 ( .A(n1032), .Z(n163) );
  BUF_X1 U128 ( .A(n1022), .Z(n188) );
  BUF_X1 U129 ( .A(n1046), .Z(n140) );
  BUF_X1 U130 ( .A(n1056), .Z(n116) );
  BUF_X1 U131 ( .A(n1027), .Z(n176) );
  BUF_X1 U132 ( .A(n1051), .Z(n128) );
  BUF_X1 U133 ( .A(n1061), .Z(n104) );
  BUF_X1 U134 ( .A(n1032), .Z(n164) );
  BUF_X1 U135 ( .A(n565), .Z(n294) );
  BUF_X1 U136 ( .A(n589), .Z(n246) );
  BUF_X1 U137 ( .A(n599), .Z(n222) );
  BUF_X1 U138 ( .A(n570), .Z(n282) );
  BUF_X1 U139 ( .A(n568), .Z(n288) );
  BUF_X1 U140 ( .A(n573), .Z(n276) );
  BUF_X1 U141 ( .A(n578), .Z(n264) );
  BUF_X1 U142 ( .A(n583), .Z(n252) );
  BUF_X1 U143 ( .A(n592), .Z(n240) );
  BUF_X1 U144 ( .A(n597), .Z(n228) );
  BUF_X1 U145 ( .A(n602), .Z(n216) );
  BUF_X1 U146 ( .A(n607), .Z(n204) );
  BUF_X1 U147 ( .A(n575), .Z(n270) );
  BUF_X1 U148 ( .A(n580), .Z(n258) );
  BUF_X1 U149 ( .A(n594), .Z(n234) );
  BUF_X1 U150 ( .A(n604), .Z(n210) );
  BUF_X1 U151 ( .A(n569), .Z(n285) );
  BUF_X1 U152 ( .A(n579), .Z(n261) );
  BUF_X1 U153 ( .A(n584), .Z(n249) );
  BUF_X1 U154 ( .A(n593), .Z(n237) );
  BUF_X1 U155 ( .A(n603), .Z(n213) );
  BUF_X1 U156 ( .A(n566), .Z(n290) );
  BUF_X1 U157 ( .A(n571), .Z(n278) );
  BUF_X1 U158 ( .A(n576), .Z(n266) );
  BUF_X1 U159 ( .A(n590), .Z(n242) );
  BUF_X1 U160 ( .A(n595), .Z(n230) );
  BUF_X1 U161 ( .A(n600), .Z(n218) );
  BUF_X1 U162 ( .A(n605), .Z(n206) );
  BUF_X1 U163 ( .A(n566), .Z(n289) );
  BUF_X1 U164 ( .A(n571), .Z(n277) );
  BUF_X1 U165 ( .A(n576), .Z(n265) );
  BUF_X1 U166 ( .A(n590), .Z(n241) );
  BUF_X1 U167 ( .A(n595), .Z(n229) );
  BUF_X1 U168 ( .A(n600), .Z(n217) );
  BUF_X1 U169 ( .A(n605), .Z(n205) );
  BUF_X1 U170 ( .A(n1022), .Z(n189) );
  BUF_X1 U171 ( .A(n1046), .Z(n141) );
  BUF_X1 U172 ( .A(n1056), .Z(n117) );
  BUF_X1 U173 ( .A(n1027), .Z(n177) );
  BUF_X1 U174 ( .A(n1051), .Z(n129) );
  BUF_X1 U175 ( .A(n1061), .Z(n105) );
  BUF_X1 U176 ( .A(n566), .Z(n291) );
  BUF_X1 U177 ( .A(n590), .Z(n243) );
  BUF_X1 U178 ( .A(n600), .Z(n219) );
  BUF_X1 U179 ( .A(n1032), .Z(n165) );
  BUF_X1 U180 ( .A(n571), .Z(n279) );
  BUF_X1 U181 ( .A(n595), .Z(n231) );
  BUF_X1 U182 ( .A(n605), .Z(n207) );
  BUF_X1 U183 ( .A(n576), .Z(n267) );
  BUF_X1 U184 ( .A(n1024), .Z(n186) );
  BUF_X1 U185 ( .A(n1029), .Z(n174) );
  BUF_X1 U186 ( .A(n1034), .Z(n162) );
  BUF_X1 U187 ( .A(n1039), .Z(n150) );
  BUF_X1 U188 ( .A(n1048), .Z(n138) );
  BUF_X1 U189 ( .A(n1053), .Z(n126) );
  BUF_X1 U190 ( .A(n1058), .Z(n114) );
  BUF_X1 U191 ( .A(n1063), .Z(n102) );
  BUF_X1 U192 ( .A(n1021), .Z(n192) );
  BUF_X1 U193 ( .A(n1045), .Z(n144) );
  BUF_X1 U194 ( .A(n1055), .Z(n120) );
  BUF_X1 U195 ( .A(n1026), .Z(n180) );
  BUF_X1 U196 ( .A(n1050), .Z(n132) );
  BUF_X1 U197 ( .A(n1060), .Z(n108) );
  BUF_X1 U198 ( .A(n1031), .Z(n168) );
  BUF_X1 U199 ( .A(n1036), .Z(n156) );
  BUF_X1 U200 ( .A(n1040), .Z(n147) );
  BUF_X1 U201 ( .A(n1025), .Z(n183) );
  BUF_X1 U202 ( .A(n1035), .Z(n159) );
  BUF_X1 U203 ( .A(n1049), .Z(n135) );
  BUF_X1 U204 ( .A(n1059), .Z(n111) );
  NAND2_X1 U205 ( .A1(n1621), .A2(n1617), .ZN(n1037) );
  NAND2_X1 U206 ( .A1(n1835), .A2(n1831), .ZN(n581) );
  BUF_X1 U207 ( .A(N347), .Z(n373) );
  BUF_X1 U208 ( .A(N347), .Z(n374) );
  BUF_X1 U209 ( .A(N348), .Z(n370) );
  BUF_X1 U210 ( .A(N348), .Z(n371) );
  BUF_X1 U211 ( .A(N350), .Z(n367) );
  BUF_X1 U212 ( .A(N350), .Z(n368) );
  BUF_X1 U213 ( .A(N351), .Z(n364) );
  BUF_X1 U214 ( .A(N351), .Z(n365) );
  BUF_X1 U215 ( .A(N352), .Z(n361) );
  BUF_X1 U216 ( .A(N352), .Z(n362) );
  BUF_X1 U217 ( .A(N354), .Z(n358) );
  BUF_X1 U218 ( .A(N354), .Z(n359) );
  BUF_X1 U219 ( .A(N355), .Z(n355) );
  BUF_X1 U220 ( .A(N355), .Z(n356) );
  BUF_X1 U221 ( .A(N356), .Z(n352) );
  BUF_X1 U222 ( .A(N356), .Z(n353) );
  BUF_X1 U223 ( .A(N358), .Z(n349) );
  BUF_X1 U224 ( .A(N358), .Z(n350) );
  BUF_X1 U225 ( .A(N359), .Z(n346) );
  BUF_X1 U226 ( .A(N359), .Z(n347) );
  BUF_X1 U227 ( .A(N360), .Z(n343) );
  BUF_X1 U228 ( .A(N360), .Z(n344) );
  BUF_X1 U229 ( .A(N362), .Z(n340) );
  BUF_X1 U230 ( .A(N362), .Z(n341) );
  BUF_X1 U231 ( .A(N363), .Z(n337) );
  BUF_X1 U232 ( .A(N363), .Z(n338) );
  BUF_X1 U233 ( .A(N364), .Z(n334) );
  BUF_X1 U234 ( .A(N364), .Z(n335) );
  BUF_X1 U235 ( .A(N366), .Z(n331) );
  BUF_X1 U236 ( .A(N366), .Z(n332) );
  BUF_X1 U237 ( .A(N367), .Z(n328) );
  BUF_X1 U238 ( .A(N367), .Z(n329) );
  BUF_X1 U239 ( .A(N368), .Z(n325) );
  BUF_X1 U240 ( .A(N368), .Z(n326) );
  BUF_X1 U241 ( .A(N370), .Z(n322) );
  BUF_X1 U242 ( .A(N370), .Z(n323) );
  BUF_X1 U243 ( .A(N371), .Z(n319) );
  BUF_X1 U244 ( .A(N371), .Z(n320) );
  BUF_X1 U245 ( .A(N372), .Z(n316) );
  BUF_X1 U246 ( .A(N372), .Z(n317) );
  BUF_X1 U247 ( .A(N343), .Z(n382) );
  BUF_X1 U248 ( .A(N343), .Z(n383) );
  BUF_X1 U249 ( .A(N344), .Z(n379) );
  BUF_X1 U250 ( .A(N344), .Z(n380) );
  BUF_X1 U251 ( .A(N346), .Z(n376) );
  BUF_X1 U252 ( .A(N346), .Z(n377) );
  BUF_X1 U253 ( .A(N374), .Z(n313) );
  BUF_X1 U254 ( .A(N374), .Z(n314) );
  BUF_X1 U255 ( .A(N375), .Z(n310) );
  BUF_X1 U256 ( .A(N375), .Z(n311) );
  BUF_X1 U257 ( .A(N376), .Z(n307) );
  BUF_X1 U258 ( .A(N376), .Z(n308) );
  BUF_X1 U259 ( .A(N378), .Z(n304) );
  BUF_X1 U260 ( .A(N378), .Z(n305) );
  BUF_X1 U261 ( .A(N379), .Z(n301) );
  BUF_X1 U262 ( .A(N379), .Z(n302) );
  BUF_X1 U263 ( .A(N380), .Z(n298) );
  BUF_X1 U264 ( .A(N380), .Z(n299) );
  BUF_X1 U265 ( .A(N382), .Z(n295) );
  BUF_X1 U266 ( .A(N382), .Z(n296) );
  BUF_X1 U267 ( .A(N310), .Z(n385) );
  BUF_X1 U268 ( .A(N310), .Z(n386) );
  AND2_X1 U269 ( .A1(n1612), .A2(n1617), .ZN(n1030) );
  AND2_X1 U270 ( .A1(n1630), .A2(n1617), .ZN(n1054) );
  AND2_X1 U271 ( .A1(n1635), .A2(n1617), .ZN(n1064) );
  AND2_X1 U272 ( .A1(n1826), .A2(n1831), .ZN(n574) );
  AND2_X1 U273 ( .A1(n1844), .A2(n1831), .ZN(n598) );
  AND2_X1 U274 ( .A1(n1849), .A2(n1831), .ZN(n608) );
  BUF_X1 U275 ( .A(n422), .Z(n35) );
  BUF_X1 U276 ( .A(n421), .Z(n32) );
  BUF_X1 U277 ( .A(n420), .Z(n29) );
  BUF_X1 U278 ( .A(n419), .Z(n26) );
  BUF_X1 U279 ( .A(n418), .Z(n23) );
  BUF_X1 U280 ( .A(n417), .Z(n20) );
  BUF_X1 U281 ( .A(n416), .Z(n17) );
  BUF_X1 U282 ( .A(n415), .Z(n14) );
  BUF_X1 U283 ( .A(n414), .Z(n11) );
  BUF_X1 U284 ( .A(n413), .Z(n8) );
  BUF_X1 U285 ( .A(n412), .Z(n5) );
  BUF_X1 U286 ( .A(n411), .Z(n2) );
  BUF_X1 U287 ( .A(n422), .Z(n34) );
  BUF_X1 U288 ( .A(n421), .Z(n31) );
  BUF_X1 U289 ( .A(n420), .Z(n28) );
  BUF_X1 U290 ( .A(n419), .Z(n25) );
  BUF_X1 U291 ( .A(n418), .Z(n22) );
  BUF_X1 U292 ( .A(n417), .Z(n19) );
  BUF_X1 U293 ( .A(n416), .Z(n16) );
  BUF_X1 U294 ( .A(n415), .Z(n13) );
  BUF_X1 U295 ( .A(n414), .Z(n10) );
  BUF_X1 U296 ( .A(n413), .Z(n7) );
  BUF_X1 U297 ( .A(n412), .Z(n4) );
  BUF_X1 U298 ( .A(n411), .Z(n1) );
  BUF_X1 U299 ( .A(n442), .Z(n95) );
  BUF_X1 U300 ( .A(n441), .Z(n92) );
  BUF_X1 U301 ( .A(n440), .Z(n89) );
  BUF_X1 U302 ( .A(n439), .Z(n86) );
  BUF_X1 U303 ( .A(n438), .Z(n83) );
  BUF_X1 U304 ( .A(n437), .Z(n80) );
  BUF_X1 U305 ( .A(n436), .Z(n77) );
  BUF_X1 U306 ( .A(n435), .Z(n74) );
  BUF_X1 U307 ( .A(n434), .Z(n71) );
  BUF_X1 U308 ( .A(n433), .Z(n68) );
  BUF_X1 U309 ( .A(n432), .Z(n65) );
  BUF_X1 U310 ( .A(n431), .Z(n62) );
  BUF_X1 U311 ( .A(n430), .Z(n59) );
  BUF_X1 U312 ( .A(n429), .Z(n56) );
  BUF_X1 U313 ( .A(n428), .Z(n53) );
  BUF_X1 U314 ( .A(n427), .Z(n50) );
  BUF_X1 U315 ( .A(n426), .Z(n47) );
  BUF_X1 U316 ( .A(n425), .Z(n44) );
  BUF_X1 U317 ( .A(n424), .Z(n41) );
  BUF_X1 U318 ( .A(n423), .Z(n38) );
  BUF_X1 U319 ( .A(n442), .Z(n94) );
  BUF_X1 U320 ( .A(n441), .Z(n91) );
  BUF_X1 U321 ( .A(n440), .Z(n88) );
  BUF_X1 U322 ( .A(n439), .Z(n85) );
  BUF_X1 U323 ( .A(n438), .Z(n82) );
  BUF_X1 U324 ( .A(n437), .Z(n79) );
  BUF_X1 U325 ( .A(n436), .Z(n76) );
  BUF_X1 U326 ( .A(n435), .Z(n73) );
  BUF_X1 U327 ( .A(n434), .Z(n70) );
  BUF_X1 U328 ( .A(n433), .Z(n67) );
  BUF_X1 U329 ( .A(n432), .Z(n64) );
  BUF_X1 U330 ( .A(n431), .Z(n61) );
  BUF_X1 U331 ( .A(n430), .Z(n58) );
  BUF_X1 U332 ( .A(n429), .Z(n55) );
  BUF_X1 U333 ( .A(n428), .Z(n52) );
  BUF_X1 U334 ( .A(n427), .Z(n49) );
  BUF_X1 U335 ( .A(n426), .Z(n46) );
  BUF_X1 U336 ( .A(n425), .Z(n43) );
  BUF_X1 U337 ( .A(n424), .Z(n40) );
  BUF_X1 U338 ( .A(n423), .Z(n37) );
  BUF_X1 U339 ( .A(N347), .Z(n375) );
  BUF_X1 U340 ( .A(N348), .Z(n372) );
  BUF_X1 U341 ( .A(N350), .Z(n369) );
  BUF_X1 U342 ( .A(N351), .Z(n366) );
  BUF_X1 U343 ( .A(N352), .Z(n363) );
  BUF_X1 U344 ( .A(N354), .Z(n360) );
  BUF_X1 U345 ( .A(N355), .Z(n357) );
  BUF_X1 U346 ( .A(N356), .Z(n354) );
  BUF_X1 U347 ( .A(N358), .Z(n351) );
  BUF_X1 U348 ( .A(N359), .Z(n348) );
  BUF_X1 U349 ( .A(N360), .Z(n345) );
  BUF_X1 U350 ( .A(N362), .Z(n342) );
  BUF_X1 U351 ( .A(N363), .Z(n339) );
  BUF_X1 U352 ( .A(N364), .Z(n336) );
  BUF_X1 U353 ( .A(N366), .Z(n333) );
  BUF_X1 U354 ( .A(N367), .Z(n330) );
  BUF_X1 U355 ( .A(N368), .Z(n327) );
  BUF_X1 U356 ( .A(N370), .Z(n324) );
  BUF_X1 U357 ( .A(N371), .Z(n321) );
  BUF_X1 U358 ( .A(N372), .Z(n318) );
  BUF_X1 U359 ( .A(N343), .Z(n384) );
  BUF_X1 U360 ( .A(N344), .Z(n381) );
  BUF_X1 U361 ( .A(N346), .Z(n378) );
  BUF_X1 U362 ( .A(N374), .Z(n315) );
  BUF_X1 U363 ( .A(N375), .Z(n312) );
  BUF_X1 U364 ( .A(N376), .Z(n309) );
  BUF_X1 U365 ( .A(N378), .Z(n306) );
  BUF_X1 U366 ( .A(N379), .Z(n303) );
  BUF_X1 U367 ( .A(N380), .Z(n300) );
  BUF_X1 U368 ( .A(N382), .Z(n297) );
  BUF_X1 U369 ( .A(N310), .Z(n387) );
  BUF_X1 U370 ( .A(n422), .Z(n36) );
  BUF_X1 U371 ( .A(n421), .Z(n33) );
  BUF_X1 U372 ( .A(n420), .Z(n30) );
  BUF_X1 U373 ( .A(n419), .Z(n27) );
  BUF_X1 U374 ( .A(n418), .Z(n24) );
  BUF_X1 U375 ( .A(n417), .Z(n21) );
  BUF_X1 U376 ( .A(n416), .Z(n18) );
  BUF_X1 U377 ( .A(n415), .Z(n15) );
  BUF_X1 U378 ( .A(n414), .Z(n12) );
  BUF_X1 U379 ( .A(n413), .Z(n9) );
  BUF_X1 U380 ( .A(n412), .Z(n6) );
  BUF_X1 U381 ( .A(n411), .Z(n3) );
  BUF_X1 U382 ( .A(n442), .Z(n96) );
  BUF_X1 U383 ( .A(n441), .Z(n93) );
  BUF_X1 U384 ( .A(n440), .Z(n90) );
  BUF_X1 U385 ( .A(n439), .Z(n87) );
  BUF_X1 U386 ( .A(n438), .Z(n84) );
  BUF_X1 U387 ( .A(n437), .Z(n81) );
  BUF_X1 U388 ( .A(n436), .Z(n78) );
  BUF_X1 U389 ( .A(n435), .Z(n75) );
  BUF_X1 U390 ( .A(n434), .Z(n72) );
  BUF_X1 U391 ( .A(n433), .Z(n69) );
  BUF_X1 U392 ( .A(n432), .Z(n66) );
  BUF_X1 U393 ( .A(n431), .Z(n63) );
  BUF_X1 U394 ( .A(n430), .Z(n60) );
  BUF_X1 U395 ( .A(n429), .Z(n57) );
  BUF_X1 U396 ( .A(n428), .Z(n54) );
  BUF_X1 U397 ( .A(n427), .Z(n51) );
  BUF_X1 U398 ( .A(n426), .Z(n48) );
  BUF_X1 U399 ( .A(n425), .Z(n45) );
  BUF_X1 U400 ( .A(n424), .Z(n42) );
  BUF_X1 U401 ( .A(n423), .Z(n39) );
  NOR2_X1 U402 ( .A1(n408), .A2(n409), .ZN(n1617) );
  NOR2_X1 U403 ( .A1(n404), .A2(n405), .ZN(n1831) );
  NOR3_X1 U404 ( .A1(ADDR_WR[3]), .A2(ADDR_WR[4]), .A3(n1003), .ZN(n969) );
  NAND2_X1 U405 ( .A1(n1615), .A2(n1621), .ZN(n1032) );
  NAND2_X1 U406 ( .A1(n1615), .A2(n1622), .ZN(n1031) );
  NAND2_X1 U407 ( .A1(n1829), .A2(n1836), .ZN(n575) );
  NAND2_X1 U408 ( .A1(n1829), .A2(n1835), .ZN(n576) );
  BUF_X1 U409 ( .A(RST), .Z(n391) );
  NAND2_X1 U410 ( .A1(n1617), .A2(n1622), .ZN(n1036) );
  NAND2_X1 U411 ( .A1(n1831), .A2(n1836), .ZN(n580) );
  NAND2_X1 U412 ( .A1(n1612), .A2(n1615), .ZN(n1022) );
  NAND2_X1 U413 ( .A1(n1614), .A2(n1615), .ZN(n1021) );
  NAND2_X1 U414 ( .A1(n1630), .A2(n1615), .ZN(n1046) );
  NAND2_X1 U415 ( .A1(n1631), .A2(n1615), .ZN(n1045) );
  NAND2_X1 U416 ( .A1(n1635), .A2(n1615), .ZN(n1056) );
  NAND2_X1 U417 ( .A1(n1636), .A2(n1615), .ZN(n1055) );
  NAND2_X1 U418 ( .A1(n1828), .A2(n1829), .ZN(n565) );
  NAND2_X1 U419 ( .A1(n1826), .A2(n1829), .ZN(n566) );
  NAND2_X1 U420 ( .A1(n1845), .A2(n1829), .ZN(n589) );
  NAND2_X1 U421 ( .A1(n1844), .A2(n1829), .ZN(n590) );
  NAND2_X1 U422 ( .A1(n1850), .A2(n1829), .ZN(n599) );
  NAND2_X1 U423 ( .A1(n1849), .A2(n1829), .ZN(n600) );
  BUF_X1 U424 ( .A(RST), .Z(n396) );
  BUF_X1 U425 ( .A(RST), .Z(n395) );
  BUF_X1 U426 ( .A(RST), .Z(n394) );
  BUF_X1 U427 ( .A(RST), .Z(n393) );
  BUF_X1 U428 ( .A(RST), .Z(n392) );
  NAND2_X1 U429 ( .A1(n1612), .A2(n1618), .ZN(n1027) );
  NAND2_X1 U430 ( .A1(n1614), .A2(n1618), .ZN(n1026) );
  NAND2_X1 U431 ( .A1(n1630), .A2(n1618), .ZN(n1051) );
  NAND2_X1 U432 ( .A1(n1631), .A2(n1618), .ZN(n1050) );
  NAND2_X1 U433 ( .A1(n1635), .A2(n1618), .ZN(n1061) );
  NAND2_X1 U434 ( .A1(n1636), .A2(n1618), .ZN(n1060) );
  NAND2_X1 U435 ( .A1(n1828), .A2(n1832), .ZN(n570) );
  NAND2_X1 U436 ( .A1(n1826), .A2(n1832), .ZN(n571) );
  NAND2_X1 U437 ( .A1(n1845), .A2(n1832), .ZN(n594) );
  NAND2_X1 U438 ( .A1(n1844), .A2(n1832), .ZN(n595) );
  NAND2_X1 U439 ( .A1(n1850), .A2(n1832), .ZN(n604) );
  NAND2_X1 U440 ( .A1(n1849), .A2(n1832), .ZN(n605) );
  OAI21_X1 U441 ( .B1(n1007), .B2(n1014), .A(n390), .ZN(N347) );
  OAI21_X1 U442 ( .B1(n1006), .B2(n1014), .A(n390), .ZN(N348) );
  OAI21_X1 U443 ( .B1(n1005), .B2(n1014), .A(n390), .ZN(N350) );
  OAI21_X1 U444 ( .B1(n1003), .B2(n1014), .A(n390), .ZN(N351) );
  OAI21_X1 U445 ( .B1(n1011), .B2(n1013), .A(n390), .ZN(N352) );
  OAI21_X1 U446 ( .B1(n1010), .B2(n1013), .A(n390), .ZN(N354) );
  OAI21_X1 U447 ( .B1(n1009), .B2(n1013), .A(n390), .ZN(N355) );
  OAI21_X1 U448 ( .B1(n1008), .B2(n1013), .A(n390), .ZN(N356) );
  OAI21_X1 U449 ( .B1(n1007), .B2(n1013), .A(n390), .ZN(N358) );
  OAI21_X1 U450 ( .B1(n1006), .B2(n1013), .A(n390), .ZN(N359) );
  OAI21_X1 U451 ( .B1(n1005), .B2(n1013), .A(n390), .ZN(N360) );
  OAI21_X1 U452 ( .B1(n1003), .B2(n1013), .A(n390), .ZN(N362) );
  OAI21_X1 U453 ( .B1(n1011), .B2(n1012), .A(n390), .ZN(N363) );
  OAI21_X1 U454 ( .B1(n1010), .B2(n1012), .A(n388), .ZN(N364) );
  OAI21_X1 U455 ( .B1(n1009), .B2(n1012), .A(n389), .ZN(N366) );
  OAI21_X1 U456 ( .B1(n1008), .B2(n1012), .A(n390), .ZN(N367) );
  OAI21_X1 U457 ( .B1(n1007), .B2(n1012), .A(n388), .ZN(N368) );
  OAI21_X1 U458 ( .B1(n1006), .B2(n1012), .A(n389), .ZN(N370) );
  OAI21_X1 U459 ( .B1(n1005), .B2(n1012), .A(n390), .ZN(N371) );
  OAI21_X1 U460 ( .B1(n1003), .B2(n1012), .A(n388), .ZN(N372) );
  OAI21_X1 U461 ( .B1(n1010), .B2(n1014), .A(n389), .ZN(N343) );
  OAI21_X1 U462 ( .B1(n1009), .B2(n1014), .A(n389), .ZN(N344) );
  OAI21_X1 U463 ( .B1(n1008), .B2(n1014), .A(n389), .ZN(N346) );
  AND2_X1 U464 ( .A1(n1624), .A2(n410), .ZN(n1621) );
  AND2_X1 U465 ( .A1(n1838), .A2(n406), .ZN(n1835) );
  AND2_X1 U466 ( .A1(n1633), .A2(n410), .ZN(n1630) );
  AND2_X1 U467 ( .A1(n1638), .A2(n410), .ZN(n1635) );
  AND2_X1 U468 ( .A1(n1847), .A2(n406), .ZN(n1844) );
  AND2_X1 U469 ( .A1(n1852), .A2(n406), .ZN(n1849) );
  AND2_X1 U470 ( .A1(n1619), .A2(n410), .ZN(n1612) );
  AND2_X1 U471 ( .A1(n1833), .A2(n406), .ZN(n1826) );
  BUF_X1 U472 ( .A(n1002), .Z(n193) );
  BUF_X1 U473 ( .A(n1002), .Z(n194) );
  AND2_X1 U474 ( .A1(n1618), .A2(n1622), .ZN(n1039) );
  AND2_X1 U475 ( .A1(n1618), .A2(n1621), .ZN(n1040) );
  AND2_X1 U476 ( .A1(n1832), .A2(n1836), .ZN(n583) );
  AND2_X1 U477 ( .A1(n1832), .A2(n1835), .ZN(n584) );
  OAI21_X1 U478 ( .B1(n1004), .B2(n1011), .A(n389), .ZN(N374) );
  OAI21_X1 U479 ( .B1(n1004), .B2(n1010), .A(n390), .ZN(N375) );
  OAI21_X1 U480 ( .B1(n1004), .B2(n1009), .A(n388), .ZN(N376) );
  OAI21_X1 U481 ( .B1(n1004), .B2(n1008), .A(n389), .ZN(N378) );
  OAI21_X1 U482 ( .B1(n1004), .B2(n1007), .A(n390), .ZN(N379) );
  OAI21_X1 U483 ( .B1(n1004), .B2(n1006), .A(n388), .ZN(N380) );
  OAI21_X1 U484 ( .B1(n1004), .B2(n1005), .A(n389), .ZN(N382) );
  AND2_X1 U485 ( .A1(n1613), .A2(n1622), .ZN(n1034) );
  AND2_X1 U486 ( .A1(n1613), .A2(n1621), .ZN(n1035) );
  AND2_X1 U487 ( .A1(n1827), .A2(n1836), .ZN(n578) );
  AND2_X1 U488 ( .A1(n1827), .A2(n1835), .ZN(n579) );
  AND2_X1 U489 ( .A1(n1614), .A2(n1617), .ZN(n1029) );
  AND2_X1 U490 ( .A1(n1631), .A2(n1617), .ZN(n1053) );
  AND2_X1 U491 ( .A1(n1636), .A2(n1617), .ZN(n1063) );
  AND2_X1 U492 ( .A1(n1828), .A2(n1831), .ZN(n573) );
  AND2_X1 U493 ( .A1(n1845), .A2(n1831), .ZN(n597) );
  AND2_X1 U494 ( .A1(n1850), .A2(n1831), .ZN(n607) );
  BUF_X1 U495 ( .A(n1002), .Z(n195) );
  AND2_X1 U496 ( .A1(n1614), .A2(n1613), .ZN(n1024) );
  AND2_X1 U497 ( .A1(n1612), .A2(n1613), .ZN(n1025) );
  AND2_X1 U498 ( .A1(n1631), .A2(n1613), .ZN(n1048) );
  AND2_X1 U499 ( .A1(n1630), .A2(n1613), .ZN(n1049) );
  AND2_X1 U500 ( .A1(n1636), .A2(n1613), .ZN(n1058) );
  AND2_X1 U501 ( .A1(n1635), .A2(n1613), .ZN(n1059) );
  AND2_X1 U502 ( .A1(n1828), .A2(n1827), .ZN(n568) );
  AND2_X1 U503 ( .A1(n1826), .A2(n1827), .ZN(n569) );
  AND2_X1 U504 ( .A1(n1845), .A2(n1827), .ZN(n592) );
  AND2_X1 U505 ( .A1(n1844), .A2(n1827), .ZN(n593) );
  AND2_X1 U506 ( .A1(n1850), .A2(n1827), .ZN(n602) );
  AND2_X1 U507 ( .A1(n1849), .A2(n1827), .ZN(n603) );
  OAI21_X1 U508 ( .B1(n1011), .B2(n1014), .A(n388), .ZN(N310) );
  NOR2_X1 U509 ( .A1(n198), .A2(n1001), .ZN(N384) );
  NOR2_X1 U510 ( .A1(n198), .A2(n1000), .ZN(N385) );
  NOR2_X1 U511 ( .A1(n198), .A2(n999), .ZN(N386) );
  NOR2_X1 U512 ( .A1(n198), .A2(n998), .ZN(N387) );
  NOR2_X1 U513 ( .A1(n198), .A2(n997), .ZN(N388) );
  NOR2_X1 U514 ( .A1(n198), .A2(n996), .ZN(N389) );
  NOR2_X1 U515 ( .A1(n198), .A2(n995), .ZN(N390) );
  NOR2_X1 U516 ( .A1(n198), .A2(n994), .ZN(N391) );
  INV_X1 U517 ( .A(ADDR_WR[2]), .ZN(n400) );
  INV_X1 U518 ( .A(ADDR_WR[0]), .ZN(n402) );
  INV_X1 U519 ( .A(ADDR_WR[1]), .ZN(n401) );
  BUF_X1 U520 ( .A(RST), .Z(n397) );
  INV_X1 U521 ( .A(n981), .ZN(n422) );
  INV_X1 U522 ( .A(n980), .ZN(n421) );
  INV_X1 U523 ( .A(n979), .ZN(n420) );
  INV_X1 U524 ( .A(n978), .ZN(n419) );
  INV_X1 U525 ( .A(n977), .ZN(n418) );
  INV_X1 U526 ( .A(n976), .ZN(n417) );
  INV_X1 U527 ( .A(n975), .ZN(n416) );
  INV_X1 U528 ( .A(n974), .ZN(n415) );
  INV_X1 U529 ( .A(n973), .ZN(n414) );
  INV_X1 U530 ( .A(n972), .ZN(n413) );
  INV_X1 U531 ( .A(n971), .ZN(n412) );
  INV_X1 U532 ( .A(n970), .ZN(n411) );
  NAND2_X1 U533 ( .A1(n1245), .A2(n1246), .ZN(N196) );
  NOR4_X1 U534 ( .A1(n1255), .A2(n1256), .A3(n1257), .A4(n1258), .ZN(n1245) );
  NOR4_X1 U535 ( .A1(n1247), .A2(n1248), .A3(n1249), .A4(n1250), .ZN(n1246) );
  OAI221_X1 U536 ( .B1(n1981), .B2(n106), .C1(n1949), .C2(n104), .A(n1262), 
        .ZN(n1255) );
  NAND2_X1 U537 ( .A1(n1263), .A2(n1264), .ZN(N195) );
  NOR4_X1 U538 ( .A1(n1273), .A2(n1274), .A3(n1275), .A4(n1276), .ZN(n1263) );
  NOR4_X1 U539 ( .A1(n1265), .A2(n1266), .A3(n1267), .A4(n1268), .ZN(n1264) );
  OAI221_X1 U540 ( .B1(n1980), .B2(n107), .C1(n1948), .C2(n104), .A(n1280), 
        .ZN(n1273) );
  NAND2_X1 U541 ( .A1(n1281), .A2(n1282), .ZN(N194) );
  NOR4_X1 U542 ( .A1(n1291), .A2(n1292), .A3(n1293), .A4(n1294), .ZN(n1281) );
  NOR4_X1 U543 ( .A1(n1283), .A2(n1284), .A3(n1285), .A4(n1286), .ZN(n1282) );
  OAI221_X1 U544 ( .B1(n1979), .B2(n107), .C1(n1947), .C2(n104), .A(n1298), 
        .ZN(n1291) );
  NAND2_X1 U545 ( .A1(n1299), .A2(n1300), .ZN(N193) );
  NOR4_X1 U546 ( .A1(n1309), .A2(n1310), .A3(n1311), .A4(n1312), .ZN(n1299) );
  NOR4_X1 U547 ( .A1(n1301), .A2(n1302), .A3(n1303), .A4(n1304), .ZN(n1300) );
  OAI221_X1 U548 ( .B1(n1978), .B2(n107), .C1(n1946), .C2(n104), .A(n1316), 
        .ZN(n1309) );
  NAND2_X1 U549 ( .A1(n1317), .A2(n1318), .ZN(N192) );
  NOR4_X1 U550 ( .A1(n1327), .A2(n1328), .A3(n1329), .A4(n1330), .ZN(n1317) );
  NOR4_X1 U551 ( .A1(n1319), .A2(n1320), .A3(n1321), .A4(n1322), .ZN(n1318) );
  OAI221_X1 U552 ( .B1(n1977), .B2(n107), .C1(n1945), .C2(n104), .A(n1334), 
        .ZN(n1327) );
  NAND2_X1 U553 ( .A1(n1335), .A2(n1336), .ZN(N191) );
  NOR4_X1 U554 ( .A1(n1345), .A2(n1346), .A3(n1347), .A4(n1348), .ZN(n1335) );
  NOR4_X1 U555 ( .A1(n1337), .A2(n1338), .A3(n1339), .A4(n1340), .ZN(n1336) );
  OAI221_X1 U556 ( .B1(n1976), .B2(n107), .C1(n1944), .C2(n104), .A(n1352), 
        .ZN(n1345) );
  NAND2_X1 U557 ( .A1(n1353), .A2(n1354), .ZN(N190) );
  NOR4_X1 U558 ( .A1(n1363), .A2(n1364), .A3(n1365), .A4(n1366), .ZN(n1353) );
  NOR4_X1 U559 ( .A1(n1355), .A2(n1356), .A3(n1357), .A4(n1358), .ZN(n1354) );
  OAI221_X1 U560 ( .B1(n1975), .B2(n107), .C1(n1943), .C2(n104), .A(n1370), 
        .ZN(n1363) );
  NAND2_X1 U561 ( .A1(n1371), .A2(n1372), .ZN(N189) );
  NOR4_X1 U562 ( .A1(n1381), .A2(n1382), .A3(n1383), .A4(n1384), .ZN(n1371) );
  NOR4_X1 U563 ( .A1(n1373), .A2(n1374), .A3(n1375), .A4(n1376), .ZN(n1372) );
  OAI221_X1 U564 ( .B1(n1974), .B2(n107), .C1(n1942), .C2(n104), .A(n1388), 
        .ZN(n1381) );
  NAND2_X1 U565 ( .A1(n1389), .A2(n1390), .ZN(N188) );
  NOR4_X1 U566 ( .A1(n1399), .A2(n1400), .A3(n1401), .A4(n1402), .ZN(n1389) );
  NOR4_X1 U567 ( .A1(n1391), .A2(n1392), .A3(n1393), .A4(n1394), .ZN(n1390) );
  OAI221_X1 U568 ( .B1(n1973), .B2(n107), .C1(n1941), .C2(n104), .A(n1406), 
        .ZN(n1399) );
  NAND2_X1 U569 ( .A1(n1407), .A2(n1408), .ZN(N187) );
  NOR4_X1 U570 ( .A1(n1417), .A2(n1418), .A3(n1419), .A4(n1420), .ZN(n1407) );
  NOR4_X1 U571 ( .A1(n1409), .A2(n1410), .A3(n1411), .A4(n1412), .ZN(n1408) );
  OAI221_X1 U572 ( .B1(n1972), .B2(n107), .C1(n1940), .C2(n103), .A(n1424), 
        .ZN(n1417) );
  NAND2_X1 U573 ( .A1(n1425), .A2(n1426), .ZN(N186) );
  NOR4_X1 U574 ( .A1(n1435), .A2(n1436), .A3(n1437), .A4(n1438), .ZN(n1425) );
  NOR4_X1 U575 ( .A1(n1427), .A2(n1428), .A3(n1429), .A4(n1430), .ZN(n1426) );
  OAI221_X1 U576 ( .B1(n1971), .B2(n107), .C1(n1939), .C2(n103), .A(n1442), 
        .ZN(n1435) );
  NAND2_X1 U577 ( .A1(n1443), .A2(n1444), .ZN(N185) );
  NOR4_X1 U578 ( .A1(n1453), .A2(n1454), .A3(n1455), .A4(n1456), .ZN(n1443) );
  NOR4_X1 U579 ( .A1(n1445), .A2(n1446), .A3(n1447), .A4(n1448), .ZN(n1444) );
  OAI221_X1 U580 ( .B1(n1970), .B2(n107), .C1(n1938), .C2(n103), .A(n1460), 
        .ZN(n1453) );
  NAND2_X1 U581 ( .A1(n1461), .A2(n1462), .ZN(N184) );
  NOR4_X1 U582 ( .A1(n1471), .A2(n1472), .A3(n1473), .A4(n1474), .ZN(n1461) );
  NOR4_X1 U583 ( .A1(n1463), .A2(n1464), .A3(n1465), .A4(n1466), .ZN(n1462) );
  OAI221_X1 U584 ( .B1(n1969), .B2(n107), .C1(n1937), .C2(n103), .A(n1478), 
        .ZN(n1471) );
  NAND2_X1 U585 ( .A1(n1479), .A2(n1480), .ZN(N183) );
  NOR4_X1 U586 ( .A1(n1489), .A2(n1490), .A3(n1491), .A4(n1492), .ZN(n1479) );
  NOR4_X1 U587 ( .A1(n1481), .A2(n1482), .A3(n1483), .A4(n1484), .ZN(n1480) );
  OAI221_X1 U588 ( .B1(n1968), .B2(n107), .C1(n1936), .C2(n103), .A(n1496), 
        .ZN(n1489) );
  NAND2_X1 U589 ( .A1(n1497), .A2(n1498), .ZN(N182) );
  NOR4_X1 U590 ( .A1(n1507), .A2(n1508), .A3(n1509), .A4(n1510), .ZN(n1497) );
  NOR4_X1 U591 ( .A1(n1499), .A2(n1500), .A3(n1501), .A4(n1502), .ZN(n1498) );
  OAI221_X1 U592 ( .B1(n1967), .B2(n108), .C1(n1935), .C2(n103), .A(n1514), 
        .ZN(n1507) );
  NAND2_X1 U593 ( .A1(n1515), .A2(n1516), .ZN(N181) );
  NOR4_X1 U594 ( .A1(n1525), .A2(n1526), .A3(n1527), .A4(n1528), .ZN(n1515) );
  NOR4_X1 U595 ( .A1(n1517), .A2(n1518), .A3(n1519), .A4(n1520), .ZN(n1516) );
  OAI221_X1 U596 ( .B1(n1966), .B2(n108), .C1(n1934), .C2(n103), .A(n1532), 
        .ZN(n1525) );
  NAND2_X1 U597 ( .A1(n1533), .A2(n1534), .ZN(N180) );
  NOR4_X1 U598 ( .A1(n1543), .A2(n1544), .A3(n1545), .A4(n1546), .ZN(n1533) );
  NOR4_X1 U599 ( .A1(n1535), .A2(n1536), .A3(n1537), .A4(n1538), .ZN(n1534) );
  OAI221_X1 U600 ( .B1(n1965), .B2(n108), .C1(n1933), .C2(n103), .A(n1550), 
        .ZN(n1543) );
  NAND2_X1 U601 ( .A1(n1551), .A2(n1552), .ZN(N179) );
  NOR4_X1 U602 ( .A1(n1561), .A2(n1562), .A3(n1563), .A4(n1564), .ZN(n1551) );
  NOR4_X1 U603 ( .A1(n1553), .A2(n1554), .A3(n1555), .A4(n1556), .ZN(n1552) );
  OAI221_X1 U604 ( .B1(n1964), .B2(n108), .C1(n1932), .C2(n103), .A(n1568), 
        .ZN(n1561) );
  NAND2_X1 U605 ( .A1(n1569), .A2(n1570), .ZN(N178) );
  NOR4_X1 U606 ( .A1(n1579), .A2(n1580), .A3(n1581), .A4(n1582), .ZN(n1569) );
  NOR4_X1 U607 ( .A1(n1571), .A2(n1572), .A3(n1573), .A4(n1574), .ZN(n1570) );
  OAI221_X1 U608 ( .B1(n1963), .B2(n108), .C1(n1931), .C2(n103), .A(n1586), 
        .ZN(n1579) );
  NAND2_X1 U609 ( .A1(n1587), .A2(n1588), .ZN(N177) );
  NOR4_X1 U610 ( .A1(n1597), .A2(n1598), .A3(n1599), .A4(n1600), .ZN(n1587) );
  NOR4_X1 U611 ( .A1(n1589), .A2(n1590), .A3(n1591), .A4(n1592), .ZN(n1588) );
  OAI221_X1 U612 ( .B1(n1962), .B2(n108), .C1(n1930), .C2(n103), .A(n1604), 
        .ZN(n1597) );
  NAND2_X1 U613 ( .A1(n1605), .A2(n1606), .ZN(N176) );
  NOR4_X1 U614 ( .A1(n1625), .A2(n1626), .A3(n1627), .A4(n1628), .ZN(n1605) );
  NOR4_X1 U615 ( .A1(n1607), .A2(n1608), .A3(n1609), .A4(n1610), .ZN(n1606) );
  OAI221_X1 U616 ( .B1(n1961), .B2(n108), .C1(n1929), .C2(n103), .A(n1637), 
        .ZN(n1625) );
  NAND2_X1 U617 ( .A1(n1639), .A2(n1640), .ZN(N110) );
  NOR4_X1 U618 ( .A1(n1649), .A2(n1650), .A3(n1651), .A4(n1652), .ZN(n1639) );
  NOR4_X1 U619 ( .A1(n1641), .A2(n1642), .A3(n1643), .A4(n1644), .ZN(n1640) );
  OAI221_X1 U620 ( .B1(n208), .B2(n1992), .C1(n205), .C2(n1960), .A(n1656), 
        .ZN(n1649) );
  NAND2_X1 U621 ( .A1(n1015), .A2(n1016), .ZN(N207) );
  NOR4_X1 U622 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1015) );
  NOR4_X1 U623 ( .A1(n1017), .A2(n1018), .A3(n1019), .A4(n1020), .ZN(n1016) );
  OAI221_X1 U624 ( .B1(n106), .B2(n1992), .C1(n105), .C2(n1960), .A(n1062), 
        .ZN(n1041) );
  NAND2_X1 U625 ( .A1(n1657), .A2(n1658), .ZN(N109) );
  NOR4_X1 U626 ( .A1(n1667), .A2(n1668), .A3(n1669), .A4(n1670), .ZN(n1657) );
  NOR4_X1 U627 ( .A1(n1659), .A2(n1660), .A3(n1661), .A4(n1662), .ZN(n1658) );
  OAI221_X1 U628 ( .B1(n208), .B2(n1991), .C1(n205), .C2(n1959), .A(n1674), 
        .ZN(n1667) );
  NAND2_X1 U629 ( .A1(n1065), .A2(n1066), .ZN(N206) );
  NOR4_X1 U630 ( .A1(n1075), .A2(n1076), .A3(n1077), .A4(n1078), .ZN(n1065) );
  NOR4_X1 U631 ( .A1(n1067), .A2(n1068), .A3(n1069), .A4(n1070), .ZN(n1066) );
  OAI221_X1 U632 ( .B1(n106), .B2(n1991), .C1(n105), .C2(n1959), .A(n1082), 
        .ZN(n1075) );
  NAND2_X1 U633 ( .A1(n1675), .A2(n1676), .ZN(N108) );
  NOR4_X1 U634 ( .A1(n1685), .A2(n1686), .A3(n1687), .A4(n1688), .ZN(n1675) );
  NOR4_X1 U635 ( .A1(n1677), .A2(n1678), .A3(n1679), .A4(n1680), .ZN(n1676) );
  OAI221_X1 U636 ( .B1(n208), .B2(n1990), .C1(n205), .C2(n1958), .A(n1692), 
        .ZN(n1685) );
  NAND2_X1 U637 ( .A1(n1083), .A2(n1084), .ZN(N205) );
  NOR4_X1 U638 ( .A1(n1093), .A2(n1094), .A3(n1095), .A4(n1096), .ZN(n1083) );
  NOR4_X1 U639 ( .A1(n1085), .A2(n1086), .A3(n1087), .A4(n1088), .ZN(n1084) );
  OAI221_X1 U640 ( .B1(n106), .B2(n1990), .C1(n105), .C2(n1958), .A(n1100), 
        .ZN(n1093) );
  NAND2_X1 U641 ( .A1(n1693), .A2(n1694), .ZN(N107) );
  NOR4_X1 U642 ( .A1(n1703), .A2(n1704), .A3(n1705), .A4(n1706), .ZN(n1693) );
  NOR4_X1 U643 ( .A1(n1695), .A2(n1696), .A3(n1697), .A4(n1698), .ZN(n1694) );
  OAI221_X1 U644 ( .B1(n208), .B2(n1989), .C1(n205), .C2(n1957), .A(n1710), 
        .ZN(n1703) );
  NAND2_X1 U645 ( .A1(n1101), .A2(n1102), .ZN(N204) );
  NOR4_X1 U646 ( .A1(n1111), .A2(n1112), .A3(n1113), .A4(n1114), .ZN(n1101) );
  NOR4_X1 U647 ( .A1(n1103), .A2(n1104), .A3(n1105), .A4(n1106), .ZN(n1102) );
  OAI221_X1 U648 ( .B1(n106), .B2(n1989), .C1(n105), .C2(n1957), .A(n1118), 
        .ZN(n1111) );
  NAND2_X1 U649 ( .A1(n1711), .A2(n1712), .ZN(N106) );
  NOR4_X1 U650 ( .A1(n1721), .A2(n1722), .A3(n1723), .A4(n1724), .ZN(n1711) );
  NOR4_X1 U651 ( .A1(n1713), .A2(n1714), .A3(n1715), .A4(n1716), .ZN(n1712) );
  OAI221_X1 U652 ( .B1(n208), .B2(n1988), .C1(n205), .C2(n1956), .A(n1728), 
        .ZN(n1721) );
  NAND2_X1 U653 ( .A1(n1119), .A2(n1120), .ZN(N203) );
  NOR4_X1 U654 ( .A1(n1129), .A2(n1130), .A3(n1131), .A4(n1132), .ZN(n1119) );
  NOR4_X1 U655 ( .A1(n1121), .A2(n1122), .A3(n1123), .A4(n1124), .ZN(n1120) );
  OAI221_X1 U656 ( .B1(n106), .B2(n1988), .C1(n105), .C2(n1956), .A(n1136), 
        .ZN(n1129) );
  NAND2_X1 U657 ( .A1(n1729), .A2(n1730), .ZN(N105) );
  NOR4_X1 U658 ( .A1(n1739), .A2(n1740), .A3(n1741), .A4(n1742), .ZN(n1729) );
  NOR4_X1 U659 ( .A1(n1731), .A2(n1732), .A3(n1733), .A4(n1734), .ZN(n1730) );
  OAI221_X1 U660 ( .B1(n208), .B2(n1987), .C1(n205), .C2(n1955), .A(n1746), 
        .ZN(n1739) );
  NAND2_X1 U661 ( .A1(n1137), .A2(n1138), .ZN(N202) );
  NOR4_X1 U662 ( .A1(n1147), .A2(n1148), .A3(n1149), .A4(n1150), .ZN(n1137) );
  NOR4_X1 U663 ( .A1(n1139), .A2(n1140), .A3(n1141), .A4(n1142), .ZN(n1138) );
  OAI221_X1 U664 ( .B1(n106), .B2(n1987), .C1(n105), .C2(n1955), .A(n1154), 
        .ZN(n1147) );
  NAND2_X1 U665 ( .A1(n1747), .A2(n1748), .ZN(N104) );
  NOR4_X1 U666 ( .A1(n1757), .A2(n1758), .A3(n1759), .A4(n1760), .ZN(n1747) );
  NOR4_X1 U667 ( .A1(n1749), .A2(n1750), .A3(n1751), .A4(n1752), .ZN(n1748) );
  OAI221_X1 U668 ( .B1(n208), .B2(n1986), .C1(n205), .C2(n1954), .A(n1764), 
        .ZN(n1757) );
  NAND2_X1 U669 ( .A1(n1155), .A2(n1156), .ZN(N201) );
  NOR4_X1 U670 ( .A1(n1165), .A2(n1166), .A3(n1167), .A4(n1168), .ZN(n1155) );
  NOR4_X1 U671 ( .A1(n1157), .A2(n1158), .A3(n1159), .A4(n1160), .ZN(n1156) );
  OAI221_X1 U672 ( .B1(n106), .B2(n1986), .C1(n105), .C2(n1954), .A(n1172), 
        .ZN(n1165) );
  NAND2_X1 U673 ( .A1(n1765), .A2(n1766), .ZN(N103) );
  NOR4_X1 U674 ( .A1(n1775), .A2(n1776), .A3(n1777), .A4(n1778), .ZN(n1765) );
  NOR4_X1 U675 ( .A1(n1767), .A2(n1768), .A3(n1769), .A4(n1770), .ZN(n1766) );
  OAI221_X1 U676 ( .B1(n208), .B2(n1985), .C1(n205), .C2(n1953), .A(n1782), 
        .ZN(n1775) );
  NAND2_X1 U677 ( .A1(n1173), .A2(n1174), .ZN(N200) );
  NOR4_X1 U678 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1173) );
  NOR4_X1 U679 ( .A1(n1175), .A2(n1176), .A3(n1177), .A4(n1178), .ZN(n1174) );
  OAI221_X1 U680 ( .B1(n106), .B2(n1985), .C1(n105), .C2(n1953), .A(n1190), 
        .ZN(n1183) );
  NAND2_X1 U681 ( .A1(n1783), .A2(n1784), .ZN(N102) );
  NOR4_X1 U682 ( .A1(n1793), .A2(n1794), .A3(n1795), .A4(n1796), .ZN(n1783) );
  NOR4_X1 U683 ( .A1(n1785), .A2(n1786), .A3(n1787), .A4(n1788), .ZN(n1784) );
  OAI221_X1 U684 ( .B1(n208), .B2(n1984), .C1(n205), .C2(n1952), .A(n1800), 
        .ZN(n1793) );
  NAND2_X1 U685 ( .A1(n1191), .A2(n1192), .ZN(N199) );
  NOR4_X1 U686 ( .A1(n1201), .A2(n1202), .A3(n1203), .A4(n1204), .ZN(n1191) );
  NOR4_X1 U687 ( .A1(n1193), .A2(n1194), .A3(n1195), .A4(n1196), .ZN(n1192) );
  OAI221_X1 U688 ( .B1(n106), .B2(n1984), .C1(n104), .C2(n1952), .A(n1208), 
        .ZN(n1201) );
  NAND2_X1 U689 ( .A1(n1801), .A2(n1802), .ZN(N101) );
  NOR4_X1 U690 ( .A1(n1811), .A2(n1812), .A3(n1813), .A4(n1814), .ZN(n1801) );
  NOR4_X1 U691 ( .A1(n1803), .A2(n1804), .A3(n1805), .A4(n1806), .ZN(n1802) );
  OAI221_X1 U692 ( .B1(n208), .B2(n1983), .C1(n205), .C2(n1951), .A(n1818), 
        .ZN(n1811) );
  NAND2_X1 U693 ( .A1(n1209), .A2(n1210), .ZN(N198) );
  NOR4_X1 U694 ( .A1(n1219), .A2(n1220), .A3(n1221), .A4(n1222), .ZN(n1209) );
  NOR4_X1 U695 ( .A1(n1211), .A2(n1212), .A3(n1213), .A4(n1214), .ZN(n1210) );
  OAI221_X1 U696 ( .B1(n106), .B2(n1983), .C1(n104), .C2(n1951), .A(n1226), 
        .ZN(n1219) );
  NAND2_X1 U697 ( .A1(n1819), .A2(n1820), .ZN(N100) );
  NOR4_X1 U698 ( .A1(n1839), .A2(n1840), .A3(n1841), .A4(n1842), .ZN(n1819) );
  NOR4_X1 U699 ( .A1(n1821), .A2(n1822), .A3(n1823), .A4(n1824), .ZN(n1820) );
  OAI221_X1 U700 ( .B1(n208), .B2(n1982), .C1(n205), .C2(n1950), .A(n1851), 
        .ZN(n1839) );
  NAND2_X1 U701 ( .A1(n1227), .A2(n1228), .ZN(N197) );
  NOR4_X1 U702 ( .A1(n1237), .A2(n1238), .A3(n1239), .A4(n1240), .ZN(n1227) );
  NOR4_X1 U703 ( .A1(n1229), .A2(n1230), .A3(n1231), .A4(n1232), .ZN(n1228) );
  OAI221_X1 U704 ( .B1(n106), .B2(n1982), .C1(n104), .C2(n1950), .A(n1244), 
        .ZN(n1237) );
  NAND2_X1 U705 ( .A1(n559), .A2(n560), .ZN(N99) );
  NOR4_X1 U706 ( .A1(n585), .A2(n586), .A3(n587), .A4(n588), .ZN(n559) );
  NOR4_X1 U707 ( .A1(n561), .A2(n562), .A3(n563), .A4(n564), .ZN(n560) );
  OAI221_X1 U708 ( .B1(n210), .B2(n1981), .C1(n207), .C2(n1949), .A(n606), 
        .ZN(n585) );
  NAND2_X1 U709 ( .A1(n609), .A2(n610), .ZN(N98) );
  NOR4_X1 U710 ( .A1(n619), .A2(n620), .A3(n621), .A4(n622), .ZN(n609) );
  NOR4_X1 U711 ( .A1(n611), .A2(n612), .A3(n613), .A4(n614), .ZN(n610) );
  OAI221_X1 U712 ( .B1(n210), .B2(n1980), .C1(n207), .C2(n1948), .A(n626), 
        .ZN(n619) );
  NAND2_X1 U713 ( .A1(n627), .A2(n628), .ZN(N97) );
  NOR4_X1 U714 ( .A1(n637), .A2(n638), .A3(n639), .A4(n640), .ZN(n627) );
  NOR4_X1 U715 ( .A1(n629), .A2(n630), .A3(n631), .A4(n632), .ZN(n628) );
  OAI221_X1 U716 ( .B1(n210), .B2(n1979), .C1(n207), .C2(n1947), .A(n644), 
        .ZN(n637) );
  NAND2_X1 U717 ( .A1(n645), .A2(n646), .ZN(N96) );
  NOR4_X1 U718 ( .A1(n655), .A2(n656), .A3(n657), .A4(n658), .ZN(n645) );
  NOR4_X1 U719 ( .A1(n647), .A2(n648), .A3(n649), .A4(n650), .ZN(n646) );
  OAI221_X1 U720 ( .B1(n210), .B2(n1978), .C1(n207), .C2(n1946), .A(n662), 
        .ZN(n655) );
  NAND2_X1 U721 ( .A1(n663), .A2(n664), .ZN(N95) );
  NOR4_X1 U722 ( .A1(n673), .A2(n674), .A3(n675), .A4(n676), .ZN(n663) );
  NOR4_X1 U723 ( .A1(n665), .A2(n666), .A3(n667), .A4(n668), .ZN(n664) );
  OAI221_X1 U724 ( .B1(n210), .B2(n1977), .C1(n207), .C2(n1945), .A(n680), 
        .ZN(n673) );
  NAND2_X1 U725 ( .A1(n681), .A2(n682), .ZN(N94) );
  NOR4_X1 U726 ( .A1(n691), .A2(n692), .A3(n693), .A4(n694), .ZN(n681) );
  NOR4_X1 U727 ( .A1(n683), .A2(n684), .A3(n685), .A4(n686), .ZN(n682) );
  OAI221_X1 U728 ( .B1(n210), .B2(n1976), .C1(n207), .C2(n1944), .A(n698), 
        .ZN(n691) );
  NAND2_X1 U729 ( .A1(n699), .A2(n700), .ZN(N93) );
  NOR4_X1 U730 ( .A1(n709), .A2(n710), .A3(n711), .A4(n712), .ZN(n699) );
  NOR4_X1 U731 ( .A1(n701), .A2(n702), .A3(n703), .A4(n704), .ZN(n700) );
  OAI221_X1 U732 ( .B1(n210), .B2(n1975), .C1(n207), .C2(n1943), .A(n716), 
        .ZN(n709) );
  NAND2_X1 U733 ( .A1(n717), .A2(n718), .ZN(N92) );
  NOR4_X1 U734 ( .A1(n727), .A2(n728), .A3(n729), .A4(n730), .ZN(n717) );
  NOR4_X1 U735 ( .A1(n719), .A2(n720), .A3(n721), .A4(n722), .ZN(n718) );
  OAI221_X1 U736 ( .B1(n210), .B2(n1974), .C1(n207), .C2(n1942), .A(n734), 
        .ZN(n727) );
  NAND2_X1 U737 ( .A1(n735), .A2(n736), .ZN(N91) );
  NOR4_X1 U738 ( .A1(n745), .A2(n746), .A3(n747), .A4(n748), .ZN(n735) );
  NOR4_X1 U739 ( .A1(n737), .A2(n738), .A3(n739), .A4(n740), .ZN(n736) );
  OAI221_X1 U740 ( .B1(n209), .B2(n1973), .C1(n206), .C2(n1941), .A(n752), 
        .ZN(n745) );
  NAND2_X1 U741 ( .A1(n753), .A2(n754), .ZN(N90) );
  NOR4_X1 U742 ( .A1(n763), .A2(n764), .A3(n765), .A4(n766), .ZN(n753) );
  NOR4_X1 U743 ( .A1(n755), .A2(n756), .A3(n757), .A4(n758), .ZN(n754) );
  OAI221_X1 U744 ( .B1(n209), .B2(n1972), .C1(n206), .C2(n1940), .A(n770), 
        .ZN(n763) );
  NAND2_X1 U745 ( .A1(n771), .A2(n772), .ZN(N89) );
  NOR4_X1 U746 ( .A1(n781), .A2(n782), .A3(n783), .A4(n784), .ZN(n771) );
  NOR4_X1 U747 ( .A1(n773), .A2(n774), .A3(n775), .A4(n776), .ZN(n772) );
  OAI221_X1 U748 ( .B1(n209), .B2(n1971), .C1(n206), .C2(n1939), .A(n788), 
        .ZN(n781) );
  NAND2_X1 U749 ( .A1(n789), .A2(n790), .ZN(N88) );
  NOR4_X1 U750 ( .A1(n799), .A2(n800), .A3(n801), .A4(n802), .ZN(n789) );
  NOR4_X1 U751 ( .A1(n791), .A2(n792), .A3(n793), .A4(n794), .ZN(n790) );
  OAI221_X1 U752 ( .B1(n209), .B2(n1970), .C1(n206), .C2(n1938), .A(n806), 
        .ZN(n799) );
  NAND2_X1 U753 ( .A1(n807), .A2(n808), .ZN(N87) );
  NOR4_X1 U754 ( .A1(n817), .A2(n818), .A3(n819), .A4(n820), .ZN(n807) );
  NOR4_X1 U755 ( .A1(n809), .A2(n810), .A3(n811), .A4(n812), .ZN(n808) );
  OAI221_X1 U756 ( .B1(n209), .B2(n1969), .C1(n206), .C2(n1937), .A(n824), 
        .ZN(n817) );
  NAND2_X1 U757 ( .A1(n825), .A2(n826), .ZN(N86) );
  NOR4_X1 U758 ( .A1(n835), .A2(n836), .A3(n837), .A4(n838), .ZN(n825) );
  NOR4_X1 U759 ( .A1(n827), .A2(n828), .A3(n829), .A4(n830), .ZN(n826) );
  OAI221_X1 U760 ( .B1(n209), .B2(n1968), .C1(n206), .C2(n1936), .A(n842), 
        .ZN(n835) );
  NAND2_X1 U761 ( .A1(n843), .A2(n844), .ZN(N85) );
  NOR4_X1 U762 ( .A1(n853), .A2(n854), .A3(n855), .A4(n856), .ZN(n843) );
  NOR4_X1 U763 ( .A1(n845), .A2(n846), .A3(n847), .A4(n848), .ZN(n844) );
  OAI221_X1 U764 ( .B1(n209), .B2(n1967), .C1(n206), .C2(n1935), .A(n860), 
        .ZN(n853) );
  NAND2_X1 U765 ( .A1(n861), .A2(n862), .ZN(N84) );
  NOR4_X1 U766 ( .A1(n871), .A2(n872), .A3(n873), .A4(n874), .ZN(n861) );
  NOR4_X1 U767 ( .A1(n863), .A2(n864), .A3(n865), .A4(n866), .ZN(n862) );
  OAI221_X1 U768 ( .B1(n209), .B2(n1966), .C1(n206), .C2(n1934), .A(n878), 
        .ZN(n871) );
  NAND2_X1 U769 ( .A1(n879), .A2(n880), .ZN(N83) );
  NOR4_X1 U770 ( .A1(n889), .A2(n890), .A3(n891), .A4(n892), .ZN(n879) );
  NOR4_X1 U771 ( .A1(n881), .A2(n882), .A3(n883), .A4(n884), .ZN(n880) );
  OAI221_X1 U772 ( .B1(n209), .B2(n1965), .C1(n206), .C2(n1933), .A(n896), 
        .ZN(n889) );
  NAND2_X1 U773 ( .A1(n897), .A2(n898), .ZN(N82) );
  NOR4_X1 U774 ( .A1(n907), .A2(n908), .A3(n909), .A4(n910), .ZN(n897) );
  NOR4_X1 U775 ( .A1(n899), .A2(n900), .A3(n901), .A4(n902), .ZN(n898) );
  OAI221_X1 U776 ( .B1(n209), .B2(n1964), .C1(n206), .C2(n1932), .A(n914), 
        .ZN(n907) );
  NAND2_X1 U777 ( .A1(n915), .A2(n916), .ZN(N81) );
  NOR4_X1 U778 ( .A1(n925), .A2(n926), .A3(n927), .A4(n928), .ZN(n915) );
  NOR4_X1 U779 ( .A1(n917), .A2(n918), .A3(n919), .A4(n920), .ZN(n916) );
  OAI221_X1 U780 ( .B1(n209), .B2(n1963), .C1(n206), .C2(n1931), .A(n932), 
        .ZN(n925) );
  NAND2_X1 U781 ( .A1(n933), .A2(n934), .ZN(N80) );
  NOR4_X1 U782 ( .A1(n943), .A2(n944), .A3(n945), .A4(n946), .ZN(n933) );
  NOR4_X1 U783 ( .A1(n935), .A2(n936), .A3(n937), .A4(n938), .ZN(n934) );
  OAI221_X1 U784 ( .B1(n209), .B2(n1962), .C1(n206), .C2(n1930), .A(n950), 
        .ZN(n943) );
  NAND2_X1 U785 ( .A1(n951), .A2(n952), .ZN(N79) );
  NOR4_X1 U786 ( .A1(n961), .A2(n962), .A3(n963), .A4(n964), .ZN(n951) );
  NOR4_X1 U787 ( .A1(n953), .A2(n954), .A3(n955), .A4(n956), .ZN(n952) );
  OAI221_X1 U788 ( .B1(n208), .B2(n1961), .C1(n205), .C2(n1929), .A(n968), 
        .ZN(n961) );
  NOR2_X1 U789 ( .A1(n196), .A2(n981), .ZN(N404) );
  NOR2_X1 U790 ( .A1(n196), .A2(n980), .ZN(N405) );
  NOR2_X1 U791 ( .A1(n196), .A2(n979), .ZN(N406) );
  NOR2_X1 U792 ( .A1(n196), .A2(n978), .ZN(N407) );
  NOR2_X1 U793 ( .A1(n196), .A2(n977), .ZN(N408) );
  NOR2_X1 U794 ( .A1(n196), .A2(n976), .ZN(N409) );
  NOR2_X1 U795 ( .A1(n196), .A2(n975), .ZN(N410) );
  NOR2_X1 U796 ( .A1(n196), .A2(n974), .ZN(N411) );
  NOR2_X1 U797 ( .A1(n196), .A2(n973), .ZN(N412) );
  NOR2_X1 U798 ( .A1(n196), .A2(n972), .ZN(N413) );
  NOR2_X1 U799 ( .A1(n196), .A2(n971), .ZN(N414) );
  NOR2_X1 U800 ( .A1(n196), .A2(n970), .ZN(N415) );
  NOR2_X1 U801 ( .A1(n197), .A2(n993), .ZN(N392) );
  NOR2_X1 U802 ( .A1(n197), .A2(n992), .ZN(N393) );
  NOR2_X1 U803 ( .A1(n197), .A2(n991), .ZN(N394) );
  NOR2_X1 U804 ( .A1(n197), .A2(n990), .ZN(N395) );
  NOR2_X1 U805 ( .A1(n197), .A2(n989), .ZN(N396) );
  NOR2_X1 U806 ( .A1(n197), .A2(n988), .ZN(N397) );
  NOR2_X1 U807 ( .A1(n197), .A2(n987), .ZN(N398) );
  NOR2_X1 U808 ( .A1(n197), .A2(n986), .ZN(N399) );
  NOR2_X1 U809 ( .A1(n197), .A2(n985), .ZN(N400) );
  NOR2_X1 U810 ( .A1(n197), .A2(n984), .ZN(N401) );
  NOR2_X1 U811 ( .A1(n197), .A2(n983), .ZN(N402) );
  NOR2_X1 U812 ( .A1(n197), .A2(n982), .ZN(N403) );
  INV_X1 U813 ( .A(n993), .ZN(n434) );
  INV_X1 U814 ( .A(n992), .ZN(n433) );
  INV_X1 U815 ( .A(n991), .ZN(n432) );
  INV_X1 U816 ( .A(n990), .ZN(n431) );
  INV_X1 U817 ( .A(n989), .ZN(n430) );
  INV_X1 U818 ( .A(n988), .ZN(n429) );
  INV_X1 U819 ( .A(n987), .ZN(n428) );
  INV_X1 U820 ( .A(n986), .ZN(n427) );
  INV_X1 U821 ( .A(n985), .ZN(n426) );
  INV_X1 U822 ( .A(n984), .ZN(n425) );
  INV_X1 U823 ( .A(n983), .ZN(n424) );
  INV_X1 U824 ( .A(n982), .ZN(n423) );
  INV_X1 U825 ( .A(n1001), .ZN(n442) );
  INV_X1 U826 ( .A(n1000), .ZN(n441) );
  INV_X1 U827 ( .A(n999), .ZN(n440) );
  INV_X1 U828 ( .A(n998), .ZN(n439) );
  INV_X1 U829 ( .A(n997), .ZN(n438) );
  INV_X1 U830 ( .A(n996), .ZN(n437) );
  INV_X1 U831 ( .A(n995), .ZN(n436) );
  INV_X1 U832 ( .A(n994), .ZN(n435) );
  INV_X1 U833 ( .A(ADDR_WR[3]), .ZN(n399) );
  INV_X1 U834 ( .A(ADDR_WR[4]), .ZN(n398) );
  NOR2_X1 U835 ( .A1(n409), .A2(ADDR_RD2[2]), .ZN(n1613) );
  NOR2_X1 U836 ( .A1(n405), .A2(ADDR_RD1[2]), .ZN(n1827) );
  OAI221_X1 U837 ( .B1(n294), .B2(n2045), .C1(n291), .C2(n2013), .A(n567), 
        .ZN(n564) );
  AOI22_X1 U838 ( .A1(\REGS[19][11] ), .A2(n288), .B1(\REGS[18][11] ), .B2(
        n285), .ZN(n567) );
  OAI221_X1 U839 ( .B1(n246), .B2(n495), .C1(n243), .C2(n463), .A(n591), .ZN(
        n588) );
  AOI22_X1 U840 ( .A1(\REGS[3][11] ), .A2(n240), .B1(\REGS[2][11] ), .B2(n237), 
        .ZN(n591) );
  OAI221_X1 U841 ( .B1(n294), .B2(n2044), .C1(n291), .C2(n2012), .A(n615), 
        .ZN(n614) );
  AOI22_X1 U842 ( .A1(\REGS[19][12] ), .A2(n288), .B1(\REGS[18][12] ), .B2(
        n285), .ZN(n615) );
  OAI221_X1 U843 ( .B1(n246), .B2(n494), .C1(n243), .C2(n462), .A(n623), .ZN(
        n622) );
  AOI22_X1 U844 ( .A1(\REGS[3][12] ), .A2(n240), .B1(\REGS[2][12] ), .B2(n237), 
        .ZN(n623) );
  OAI221_X1 U845 ( .B1(n294), .B2(n2043), .C1(n291), .C2(n2011), .A(n633), 
        .ZN(n632) );
  AOI22_X1 U846 ( .A1(\REGS[19][13] ), .A2(n288), .B1(\REGS[18][13] ), .B2(
        n285), .ZN(n633) );
  OAI221_X1 U847 ( .B1(n246), .B2(n493), .C1(n243), .C2(n461), .A(n641), .ZN(
        n640) );
  AOI22_X1 U848 ( .A1(\REGS[3][13] ), .A2(n240), .B1(\REGS[2][13] ), .B2(n237), 
        .ZN(n641) );
  OAI221_X1 U849 ( .B1(n294), .B2(n2042), .C1(n291), .C2(n2010), .A(n651), 
        .ZN(n650) );
  AOI22_X1 U850 ( .A1(\REGS[19][14] ), .A2(n288), .B1(\REGS[18][14] ), .B2(
        n285), .ZN(n651) );
  OAI221_X1 U851 ( .B1(n246), .B2(n492), .C1(n243), .C2(n460), .A(n659), .ZN(
        n658) );
  AOI22_X1 U852 ( .A1(\REGS[3][14] ), .A2(n240), .B1(\REGS[2][14] ), .B2(n237), 
        .ZN(n659) );
  OAI221_X1 U853 ( .B1(n294), .B2(n2041), .C1(n291), .C2(n2009), .A(n669), 
        .ZN(n668) );
  AOI22_X1 U854 ( .A1(\REGS[19][15] ), .A2(n288), .B1(\REGS[18][15] ), .B2(
        n285), .ZN(n669) );
  OAI221_X1 U855 ( .B1(n246), .B2(n491), .C1(n243), .C2(n459), .A(n677), .ZN(
        n676) );
  AOI22_X1 U856 ( .A1(\REGS[3][15] ), .A2(n240), .B1(\REGS[2][15] ), .B2(n237), 
        .ZN(n677) );
  OAI221_X1 U857 ( .B1(n294), .B2(n2040), .C1(n291), .C2(n2008), .A(n687), 
        .ZN(n686) );
  AOI22_X1 U858 ( .A1(\REGS[19][16] ), .A2(n288), .B1(\REGS[18][16] ), .B2(
        n285), .ZN(n687) );
  OAI221_X1 U859 ( .B1(n246), .B2(n490), .C1(n243), .C2(n458), .A(n695), .ZN(
        n694) );
  AOI22_X1 U860 ( .A1(\REGS[3][16] ), .A2(n240), .B1(\REGS[2][16] ), .B2(n237), 
        .ZN(n695) );
  OAI221_X1 U861 ( .B1(n294), .B2(n2039), .C1(n291), .C2(n2007), .A(n705), 
        .ZN(n704) );
  AOI22_X1 U862 ( .A1(\REGS[19][17] ), .A2(n288), .B1(\REGS[18][17] ), .B2(
        n285), .ZN(n705) );
  OAI221_X1 U863 ( .B1(n246), .B2(n489), .C1(n243), .C2(n457), .A(n713), .ZN(
        n712) );
  AOI22_X1 U864 ( .A1(\REGS[3][17] ), .A2(n240), .B1(\REGS[2][17] ), .B2(n237), 
        .ZN(n713) );
  OAI221_X1 U865 ( .B1(n294), .B2(n2038), .C1(n291), .C2(n2006), .A(n723), 
        .ZN(n722) );
  AOI22_X1 U866 ( .A1(\REGS[19][18] ), .A2(n288), .B1(\REGS[18][18] ), .B2(
        n285), .ZN(n723) );
  OAI221_X1 U867 ( .B1(n246), .B2(n488), .C1(n243), .C2(n456), .A(n731), .ZN(
        n730) );
  AOI22_X1 U868 ( .A1(\REGS[3][18] ), .A2(n240), .B1(\REGS[2][18] ), .B2(n237), 
        .ZN(n731) );
  OAI221_X1 U869 ( .B1(n2031), .B2(n192), .C1(n1999), .C2(n187), .A(n1503), 
        .ZN(n1502) );
  AOI22_X1 U870 ( .A1(n186), .A2(\REGS[19][25] ), .B1(n183), .B2(
        \REGS[18][25] ), .ZN(n1503) );
  OAI221_X1 U871 ( .B1(n481), .B2(n144), .C1(n449), .C2(n139), .A(n1511), .ZN(
        n1510) );
  AOI22_X1 U872 ( .A1(n138), .A2(\REGS[3][25] ), .B1(n135), .B2(\REGS[2][25] ), 
        .ZN(n1511) );
  OAI221_X1 U873 ( .B1(n2030), .B2(n192), .C1(n1998), .C2(n187), .A(n1521), 
        .ZN(n1520) );
  AOI22_X1 U874 ( .A1(n186), .A2(\REGS[19][26] ), .B1(n183), .B2(
        \REGS[18][26] ), .ZN(n1521) );
  OAI221_X1 U875 ( .B1(n480), .B2(n144), .C1(n448), .C2(n139), .A(n1529), .ZN(
        n1528) );
  AOI22_X1 U876 ( .A1(n138), .A2(\REGS[3][26] ), .B1(n135), .B2(\REGS[2][26] ), 
        .ZN(n1529) );
  OAI221_X1 U877 ( .B1(n2029), .B2(n192), .C1(n1997), .C2(n187), .A(n1539), 
        .ZN(n1538) );
  AOI22_X1 U878 ( .A1(n186), .A2(\REGS[19][27] ), .B1(n183), .B2(
        \REGS[18][27] ), .ZN(n1539) );
  OAI221_X1 U879 ( .B1(n479), .B2(n144), .C1(n447), .C2(n139), .A(n1547), .ZN(
        n1546) );
  AOI22_X1 U880 ( .A1(n138), .A2(\REGS[3][27] ), .B1(n135), .B2(\REGS[2][27] ), 
        .ZN(n1547) );
  OAI221_X1 U881 ( .B1(n2028), .B2(n192), .C1(n1996), .C2(n187), .A(n1557), 
        .ZN(n1556) );
  AOI22_X1 U882 ( .A1(n186), .A2(\REGS[19][28] ), .B1(n183), .B2(
        \REGS[18][28] ), .ZN(n1557) );
  OAI221_X1 U883 ( .B1(n478), .B2(n144), .C1(n446), .C2(n139), .A(n1565), .ZN(
        n1564) );
  AOI22_X1 U884 ( .A1(n138), .A2(\REGS[3][28] ), .B1(n135), .B2(\REGS[2][28] ), 
        .ZN(n1565) );
  OAI221_X1 U885 ( .B1(n2027), .B2(n192), .C1(n1995), .C2(n187), .A(n1575), 
        .ZN(n1574) );
  AOI22_X1 U886 ( .A1(n186), .A2(\REGS[19][29] ), .B1(n183), .B2(
        \REGS[18][29] ), .ZN(n1575) );
  OAI221_X1 U887 ( .B1(n477), .B2(n144), .C1(n445), .C2(n139), .A(n1583), .ZN(
        n1582) );
  AOI22_X1 U888 ( .A1(n138), .A2(\REGS[3][29] ), .B1(n135), .B2(\REGS[2][29] ), 
        .ZN(n1583) );
  OAI221_X1 U889 ( .B1(n2026), .B2(n192), .C1(n1994), .C2(n187), .A(n1593), 
        .ZN(n1592) );
  AOI22_X1 U890 ( .A1(n186), .A2(\REGS[19][30] ), .B1(n183), .B2(
        \REGS[18][30] ), .ZN(n1593) );
  OAI221_X1 U891 ( .B1(n476), .B2(n144), .C1(n444), .C2(n139), .A(n1601), .ZN(
        n1600) );
  AOI22_X1 U892 ( .A1(n138), .A2(\REGS[3][30] ), .B1(n135), .B2(\REGS[2][30] ), 
        .ZN(n1601) );
  OAI221_X1 U893 ( .B1(n2025), .B2(n192), .C1(n1993), .C2(n187), .A(n1611), 
        .ZN(n1610) );
  AOI22_X1 U894 ( .A1(n186), .A2(\REGS[19][31] ), .B1(n183), .B2(
        \REGS[18][31] ), .ZN(n1611) );
  OAI221_X1 U895 ( .B1(n475), .B2(n144), .C1(n443), .C2(n139), .A(n1629), .ZN(
        n1628) );
  AOI22_X1 U896 ( .A1(n138), .A2(\REGS[3][31] ), .B1(n135), .B2(\REGS[2][31] ), 
        .ZN(n1629) );
  OAI221_X1 U897 ( .B1(n292), .B2(n2056), .C1(n289), .C2(n2024), .A(n1645), 
        .ZN(n1644) );
  AOI22_X1 U898 ( .A1(\REGS[19][0] ), .A2(n286), .B1(\REGS[18][0] ), .B2(n283), 
        .ZN(n1645) );
  OAI221_X1 U899 ( .B1(n244), .B2(n506), .C1(n241), .C2(n474), .A(n1653), .ZN(
        n1652) );
  AOI22_X1 U900 ( .A1(\REGS[3][0] ), .A2(n238), .B1(\REGS[2][0] ), .B2(n235), 
        .ZN(n1653) );
  OAI221_X1 U901 ( .B1(n190), .B2(n2056), .C1(n189), .C2(n2024), .A(n1023), 
        .ZN(n1020) );
  AOI22_X1 U902 ( .A1(\REGS[19][0] ), .A2(n184), .B1(\REGS[18][0] ), .B2(n181), 
        .ZN(n1023) );
  OAI221_X1 U903 ( .B1(n142), .B2(n506), .C1(n141), .C2(n474), .A(n1047), .ZN(
        n1044) );
  AOI22_X1 U904 ( .A1(\REGS[3][0] ), .A2(n136), .B1(\REGS[2][0] ), .B2(n133), 
        .ZN(n1047) );
  OAI221_X1 U905 ( .B1(n292), .B2(n2055), .C1(n289), .C2(n2023), .A(n1663), 
        .ZN(n1662) );
  AOI22_X1 U906 ( .A1(\REGS[19][1] ), .A2(n286), .B1(\REGS[18][1] ), .B2(n283), 
        .ZN(n1663) );
  OAI221_X1 U907 ( .B1(n244), .B2(n505), .C1(n241), .C2(n473), .A(n1671), .ZN(
        n1670) );
  AOI22_X1 U908 ( .A1(\REGS[3][1] ), .A2(n238), .B1(\REGS[2][1] ), .B2(n235), 
        .ZN(n1671) );
  OAI221_X1 U909 ( .B1(n190), .B2(n2055), .C1(n189), .C2(n2023), .A(n1071), 
        .ZN(n1070) );
  AOI22_X1 U910 ( .A1(\REGS[19][1] ), .A2(n184), .B1(\REGS[18][1] ), .B2(n181), 
        .ZN(n1071) );
  OAI221_X1 U911 ( .B1(n142), .B2(n505), .C1(n141), .C2(n473), .A(n1079), .ZN(
        n1078) );
  AOI22_X1 U912 ( .A1(\REGS[3][1] ), .A2(n136), .B1(\REGS[2][1] ), .B2(n133), 
        .ZN(n1079) );
  OAI221_X1 U913 ( .B1(n292), .B2(n2054), .C1(n289), .C2(n2022), .A(n1681), 
        .ZN(n1680) );
  AOI22_X1 U914 ( .A1(\REGS[19][2] ), .A2(n286), .B1(\REGS[18][2] ), .B2(n283), 
        .ZN(n1681) );
  OAI221_X1 U915 ( .B1(n244), .B2(n504), .C1(n241), .C2(n472), .A(n1689), .ZN(
        n1688) );
  AOI22_X1 U916 ( .A1(\REGS[3][2] ), .A2(n238), .B1(\REGS[2][2] ), .B2(n235), 
        .ZN(n1689) );
  OAI221_X1 U917 ( .B1(n190), .B2(n2054), .C1(n189), .C2(n2022), .A(n1089), 
        .ZN(n1088) );
  AOI22_X1 U918 ( .A1(\REGS[19][2] ), .A2(n184), .B1(\REGS[18][2] ), .B2(n181), 
        .ZN(n1089) );
  OAI221_X1 U919 ( .B1(n142), .B2(n504), .C1(n141), .C2(n472), .A(n1097), .ZN(
        n1096) );
  AOI22_X1 U920 ( .A1(\REGS[3][2] ), .A2(n136), .B1(\REGS[2][2] ), .B2(n133), 
        .ZN(n1097) );
  OAI221_X1 U921 ( .B1(n292), .B2(n2053), .C1(n289), .C2(n2021), .A(n1699), 
        .ZN(n1698) );
  AOI22_X1 U922 ( .A1(\REGS[19][3] ), .A2(n286), .B1(\REGS[18][3] ), .B2(n283), 
        .ZN(n1699) );
  OAI221_X1 U923 ( .B1(n244), .B2(n503), .C1(n241), .C2(n471), .A(n1707), .ZN(
        n1706) );
  AOI22_X1 U924 ( .A1(\REGS[3][3] ), .A2(n238), .B1(\REGS[2][3] ), .B2(n235), 
        .ZN(n1707) );
  OAI221_X1 U925 ( .B1(n190), .B2(n2053), .C1(n189), .C2(n2021), .A(n1107), 
        .ZN(n1106) );
  AOI22_X1 U926 ( .A1(\REGS[19][3] ), .A2(n184), .B1(\REGS[18][3] ), .B2(n181), 
        .ZN(n1107) );
  OAI221_X1 U927 ( .B1(n142), .B2(n503), .C1(n141), .C2(n471), .A(n1115), .ZN(
        n1114) );
  AOI22_X1 U928 ( .A1(\REGS[3][3] ), .A2(n136), .B1(\REGS[2][3] ), .B2(n133), 
        .ZN(n1115) );
  OAI221_X1 U929 ( .B1(n292), .B2(n2052), .C1(n289), .C2(n2020), .A(n1717), 
        .ZN(n1716) );
  AOI22_X1 U930 ( .A1(\REGS[19][4] ), .A2(n286), .B1(\REGS[18][4] ), .B2(n283), 
        .ZN(n1717) );
  OAI221_X1 U931 ( .B1(n244), .B2(n502), .C1(n241), .C2(n470), .A(n1725), .ZN(
        n1724) );
  AOI22_X1 U932 ( .A1(\REGS[3][4] ), .A2(n238), .B1(\REGS[2][4] ), .B2(n235), 
        .ZN(n1725) );
  OAI221_X1 U933 ( .B1(n190), .B2(n2052), .C1(n189), .C2(n2020), .A(n1125), 
        .ZN(n1124) );
  AOI22_X1 U934 ( .A1(\REGS[19][4] ), .A2(n184), .B1(\REGS[18][4] ), .B2(n181), 
        .ZN(n1125) );
  OAI221_X1 U935 ( .B1(n142), .B2(n502), .C1(n141), .C2(n470), .A(n1133), .ZN(
        n1132) );
  AOI22_X1 U936 ( .A1(\REGS[3][4] ), .A2(n136), .B1(\REGS[2][4] ), .B2(n133), 
        .ZN(n1133) );
  OAI221_X1 U937 ( .B1(n292), .B2(n2051), .C1(n289), .C2(n2019), .A(n1735), 
        .ZN(n1734) );
  AOI22_X1 U938 ( .A1(\REGS[19][5] ), .A2(n286), .B1(\REGS[18][5] ), .B2(n283), 
        .ZN(n1735) );
  OAI221_X1 U939 ( .B1(n244), .B2(n501), .C1(n241), .C2(n469), .A(n1743), .ZN(
        n1742) );
  AOI22_X1 U940 ( .A1(\REGS[3][5] ), .A2(n238), .B1(\REGS[2][5] ), .B2(n235), 
        .ZN(n1743) );
  OAI221_X1 U941 ( .B1(n190), .B2(n2051), .C1(n189), .C2(n2019), .A(n1143), 
        .ZN(n1142) );
  AOI22_X1 U942 ( .A1(\REGS[19][5] ), .A2(n184), .B1(\REGS[18][5] ), .B2(n181), 
        .ZN(n1143) );
  OAI221_X1 U943 ( .B1(n142), .B2(n501), .C1(n141), .C2(n469), .A(n1151), .ZN(
        n1150) );
  AOI22_X1 U944 ( .A1(\REGS[3][5] ), .A2(n136), .B1(\REGS[2][5] ), .B2(n133), 
        .ZN(n1151) );
  OAI221_X1 U945 ( .B1(n292), .B2(n2050), .C1(n289), .C2(n2018), .A(n1753), 
        .ZN(n1752) );
  AOI22_X1 U946 ( .A1(\REGS[19][6] ), .A2(n286), .B1(\REGS[18][6] ), .B2(n283), 
        .ZN(n1753) );
  OAI221_X1 U947 ( .B1(n244), .B2(n500), .C1(n241), .C2(n468), .A(n1761), .ZN(
        n1760) );
  AOI22_X1 U948 ( .A1(\REGS[3][6] ), .A2(n238), .B1(\REGS[2][6] ), .B2(n235), 
        .ZN(n1761) );
  OAI221_X1 U949 ( .B1(n190), .B2(n2050), .C1(n189), .C2(n2018), .A(n1161), 
        .ZN(n1160) );
  AOI22_X1 U950 ( .A1(\REGS[19][6] ), .A2(n184), .B1(\REGS[18][6] ), .B2(n181), 
        .ZN(n1161) );
  OAI221_X1 U951 ( .B1(n142), .B2(n500), .C1(n141), .C2(n468), .A(n1169), .ZN(
        n1168) );
  AOI22_X1 U952 ( .A1(\REGS[3][6] ), .A2(n136), .B1(\REGS[2][6] ), .B2(n133), 
        .ZN(n1169) );
  OAI221_X1 U953 ( .B1(n292), .B2(n2049), .C1(n289), .C2(n2017), .A(n1771), 
        .ZN(n1770) );
  AOI22_X1 U954 ( .A1(\REGS[19][7] ), .A2(n286), .B1(\REGS[18][7] ), .B2(n283), 
        .ZN(n1771) );
  OAI221_X1 U955 ( .B1(n244), .B2(n499), .C1(n241), .C2(n467), .A(n1779), .ZN(
        n1778) );
  AOI22_X1 U956 ( .A1(\REGS[3][7] ), .A2(n238), .B1(\REGS[2][7] ), .B2(n235), 
        .ZN(n1779) );
  OAI221_X1 U957 ( .B1(n190), .B2(n2049), .C1(n189), .C2(n2017), .A(n1179), 
        .ZN(n1178) );
  AOI22_X1 U958 ( .A1(\REGS[19][7] ), .A2(n184), .B1(\REGS[18][7] ), .B2(n181), 
        .ZN(n1179) );
  OAI221_X1 U959 ( .B1(n142), .B2(n499), .C1(n141), .C2(n467), .A(n1187), .ZN(
        n1186) );
  AOI22_X1 U960 ( .A1(\REGS[3][7] ), .A2(n136), .B1(\REGS[2][7] ), .B2(n133), 
        .ZN(n1187) );
  OAI221_X1 U961 ( .B1(n292), .B2(n2048), .C1(n289), .C2(n2016), .A(n1789), 
        .ZN(n1788) );
  AOI22_X1 U962 ( .A1(\REGS[19][8] ), .A2(n286), .B1(\REGS[18][8] ), .B2(n283), 
        .ZN(n1789) );
  OAI221_X1 U963 ( .B1(n244), .B2(n498), .C1(n241), .C2(n466), .A(n1797), .ZN(
        n1796) );
  AOI22_X1 U964 ( .A1(\REGS[3][8] ), .A2(n238), .B1(\REGS[2][8] ), .B2(n235), 
        .ZN(n1797) );
  OAI221_X1 U965 ( .B1(n190), .B2(n2048), .C1(n188), .C2(n2016), .A(n1197), 
        .ZN(n1196) );
  AOI22_X1 U966 ( .A1(\REGS[19][8] ), .A2(n184), .B1(\REGS[18][8] ), .B2(n181), 
        .ZN(n1197) );
  OAI221_X1 U967 ( .B1(n142), .B2(n498), .C1(n140), .C2(n466), .A(n1205), .ZN(
        n1204) );
  AOI22_X1 U968 ( .A1(\REGS[3][8] ), .A2(n136), .B1(\REGS[2][8] ), .B2(n133), 
        .ZN(n1205) );
  OAI221_X1 U969 ( .B1(n292), .B2(n2047), .C1(n289), .C2(n2015), .A(n1807), 
        .ZN(n1806) );
  AOI22_X1 U970 ( .A1(\REGS[19][9] ), .A2(n286), .B1(\REGS[18][9] ), .B2(n283), 
        .ZN(n1807) );
  OAI221_X1 U971 ( .B1(n244), .B2(n497), .C1(n241), .C2(n465), .A(n1815), .ZN(
        n1814) );
  AOI22_X1 U972 ( .A1(\REGS[3][9] ), .A2(n238), .B1(\REGS[2][9] ), .B2(n235), 
        .ZN(n1815) );
  OAI221_X1 U973 ( .B1(n190), .B2(n2047), .C1(n188), .C2(n2015), .A(n1215), 
        .ZN(n1214) );
  AOI22_X1 U974 ( .A1(\REGS[19][9] ), .A2(n184), .B1(\REGS[18][9] ), .B2(n181), 
        .ZN(n1215) );
  OAI221_X1 U975 ( .B1(n142), .B2(n497), .C1(n140), .C2(n465), .A(n1223), .ZN(
        n1222) );
  AOI22_X1 U976 ( .A1(\REGS[3][9] ), .A2(n136), .B1(\REGS[2][9] ), .B2(n133), 
        .ZN(n1223) );
  OAI221_X1 U977 ( .B1(n292), .B2(n2046), .C1(n289), .C2(n2014), .A(n1825), 
        .ZN(n1824) );
  AOI22_X1 U978 ( .A1(\REGS[19][10] ), .A2(n286), .B1(\REGS[18][10] ), .B2(
        n283), .ZN(n1825) );
  OAI221_X1 U979 ( .B1(n244), .B2(n496), .C1(n241), .C2(n464), .A(n1843), .ZN(
        n1842) );
  AOI22_X1 U980 ( .A1(\REGS[3][10] ), .A2(n238), .B1(\REGS[2][10] ), .B2(n235), 
        .ZN(n1843) );
  OAI221_X1 U981 ( .B1(n190), .B2(n2046), .C1(n188), .C2(n2014), .A(n1233), 
        .ZN(n1232) );
  AOI22_X1 U982 ( .A1(\REGS[19][10] ), .A2(n184), .B1(\REGS[18][10] ), .B2(
        n181), .ZN(n1233) );
  OAI221_X1 U983 ( .B1(n142), .B2(n496), .C1(n140), .C2(n464), .A(n1241), .ZN(
        n1240) );
  AOI22_X1 U984 ( .A1(\REGS[3][10] ), .A2(n136), .B1(\REGS[2][10] ), .B2(n133), 
        .ZN(n1241) );
  OAI221_X1 U985 ( .B1(n2045), .B2(n190), .C1(n2013), .C2(n188), .A(n1251), 
        .ZN(n1250) );
  AOI22_X1 U986 ( .A1(n184), .A2(\REGS[19][11] ), .B1(n181), .B2(
        \REGS[18][11] ), .ZN(n1251) );
  OAI221_X1 U987 ( .B1(n495), .B2(n142), .C1(n463), .C2(n140), .A(n1259), .ZN(
        n1258) );
  AOI22_X1 U988 ( .A1(n136), .A2(\REGS[3][11] ), .B1(n133), .B2(\REGS[2][11] ), 
        .ZN(n1259) );
  OAI221_X1 U989 ( .B1(n2044), .B2(n191), .C1(n2012), .C2(n188), .A(n1269), 
        .ZN(n1268) );
  AOI22_X1 U990 ( .A1(n185), .A2(\REGS[19][12] ), .B1(n182), .B2(
        \REGS[18][12] ), .ZN(n1269) );
  OAI221_X1 U991 ( .B1(n494), .B2(n143), .C1(n462), .C2(n140), .A(n1277), .ZN(
        n1276) );
  AOI22_X1 U992 ( .A1(n137), .A2(\REGS[3][12] ), .B1(n134), .B2(\REGS[2][12] ), 
        .ZN(n1277) );
  OAI221_X1 U993 ( .B1(n2043), .B2(n191), .C1(n2011), .C2(n188), .A(n1287), 
        .ZN(n1286) );
  AOI22_X1 U994 ( .A1(n185), .A2(\REGS[19][13] ), .B1(n182), .B2(
        \REGS[18][13] ), .ZN(n1287) );
  OAI221_X1 U995 ( .B1(n493), .B2(n143), .C1(n461), .C2(n140), .A(n1295), .ZN(
        n1294) );
  AOI22_X1 U996 ( .A1(n137), .A2(\REGS[3][13] ), .B1(n134), .B2(\REGS[2][13] ), 
        .ZN(n1295) );
  OAI221_X1 U997 ( .B1(n2042), .B2(n191), .C1(n2010), .C2(n188), .A(n1305), 
        .ZN(n1304) );
  AOI22_X1 U998 ( .A1(n185), .A2(\REGS[19][14] ), .B1(n182), .B2(
        \REGS[18][14] ), .ZN(n1305) );
  OAI221_X1 U999 ( .B1(n492), .B2(n143), .C1(n460), .C2(n140), .A(n1313), .ZN(
        n1312) );
  AOI22_X1 U1000 ( .A1(n137), .A2(\REGS[3][14] ), .B1(n134), .B2(\REGS[2][14] ), .ZN(n1313) );
  OAI221_X1 U1001 ( .B1(n2041), .B2(n191), .C1(n2009), .C2(n188), .A(n1323), 
        .ZN(n1322) );
  AOI22_X1 U1002 ( .A1(n185), .A2(\REGS[19][15] ), .B1(n182), .B2(
        \REGS[18][15] ), .ZN(n1323) );
  OAI221_X1 U1003 ( .B1(n491), .B2(n143), .C1(n459), .C2(n140), .A(n1331), 
        .ZN(n1330) );
  AOI22_X1 U1004 ( .A1(n137), .A2(\REGS[3][15] ), .B1(n134), .B2(\REGS[2][15] ), .ZN(n1331) );
  OAI221_X1 U1005 ( .B1(n2040), .B2(n191), .C1(n2008), .C2(n188), .A(n1341), 
        .ZN(n1340) );
  AOI22_X1 U1006 ( .A1(n185), .A2(\REGS[19][16] ), .B1(n182), .B2(
        \REGS[18][16] ), .ZN(n1341) );
  OAI221_X1 U1007 ( .B1(n490), .B2(n143), .C1(n458), .C2(n140), .A(n1349), 
        .ZN(n1348) );
  AOI22_X1 U1008 ( .A1(n137), .A2(\REGS[3][16] ), .B1(n134), .B2(\REGS[2][16] ), .ZN(n1349) );
  OAI221_X1 U1009 ( .B1(n2039), .B2(n191), .C1(n2007), .C2(n188), .A(n1359), 
        .ZN(n1358) );
  AOI22_X1 U1010 ( .A1(n185), .A2(\REGS[19][17] ), .B1(n182), .B2(
        \REGS[18][17] ), .ZN(n1359) );
  OAI221_X1 U1011 ( .B1(n489), .B2(n143), .C1(n457), .C2(n140), .A(n1367), 
        .ZN(n1366) );
  AOI22_X1 U1012 ( .A1(n137), .A2(\REGS[3][17] ), .B1(n134), .B2(\REGS[2][17] ), .ZN(n1367) );
  OAI221_X1 U1013 ( .B1(n2038), .B2(n191), .C1(n2006), .C2(n188), .A(n1377), 
        .ZN(n1376) );
  AOI22_X1 U1014 ( .A1(n185), .A2(\REGS[19][18] ), .B1(n182), .B2(
        \REGS[18][18] ), .ZN(n1377) );
  OAI221_X1 U1015 ( .B1(n488), .B2(n143), .C1(n456), .C2(n140), .A(n1385), 
        .ZN(n1384) );
  AOI22_X1 U1016 ( .A1(n137), .A2(\REGS[3][18] ), .B1(n134), .B2(\REGS[2][18] ), .ZN(n1385) );
  OAI221_X1 U1017 ( .B1(n2037), .B2(n191), .C1(n2005), .C2(n188), .A(n1395), 
        .ZN(n1394) );
  AOI22_X1 U1018 ( .A1(n185), .A2(\REGS[19][19] ), .B1(n182), .B2(
        \REGS[18][19] ), .ZN(n1395) );
  OAI221_X1 U1019 ( .B1(n487), .B2(n143), .C1(n455), .C2(n140), .A(n1403), 
        .ZN(n1402) );
  AOI22_X1 U1020 ( .A1(n137), .A2(\REGS[3][19] ), .B1(n134), .B2(\REGS[2][19] ), .ZN(n1403) );
  OAI221_X1 U1021 ( .B1(n293), .B2(n2037), .C1(n290), .C2(n2005), .A(n741), 
        .ZN(n740) );
  AOI22_X1 U1022 ( .A1(\REGS[19][19] ), .A2(n287), .B1(\REGS[18][19] ), .B2(
        n284), .ZN(n741) );
  OAI221_X1 U1023 ( .B1(n245), .B2(n487), .C1(n242), .C2(n455), .A(n749), .ZN(
        n748) );
  AOI22_X1 U1024 ( .A1(\REGS[3][19] ), .A2(n239), .B1(\REGS[2][19] ), .B2(n236), .ZN(n749) );
  OAI221_X1 U1025 ( .B1(n2036), .B2(n191), .C1(n2004), .C2(n187), .A(n1413), 
        .ZN(n1412) );
  AOI22_X1 U1026 ( .A1(n185), .A2(\REGS[19][20] ), .B1(n182), .B2(
        \REGS[18][20] ), .ZN(n1413) );
  OAI221_X1 U1027 ( .B1(n486), .B2(n143), .C1(n454), .C2(n139), .A(n1421), 
        .ZN(n1420) );
  AOI22_X1 U1028 ( .A1(n137), .A2(\REGS[3][20] ), .B1(n134), .B2(\REGS[2][20] ), .ZN(n1421) );
  OAI221_X1 U1029 ( .B1(n293), .B2(n2036), .C1(n290), .C2(n2004), .A(n759), 
        .ZN(n758) );
  AOI22_X1 U1030 ( .A1(\REGS[19][20] ), .A2(n287), .B1(\REGS[18][20] ), .B2(
        n284), .ZN(n759) );
  OAI221_X1 U1031 ( .B1(n245), .B2(n486), .C1(n242), .C2(n454), .A(n767), .ZN(
        n766) );
  AOI22_X1 U1032 ( .A1(\REGS[3][20] ), .A2(n239), .B1(\REGS[2][20] ), .B2(n236), .ZN(n767) );
  OAI221_X1 U1033 ( .B1(n2035), .B2(n191), .C1(n2003), .C2(n187), .A(n1431), 
        .ZN(n1430) );
  AOI22_X1 U1034 ( .A1(n185), .A2(\REGS[19][21] ), .B1(n182), .B2(
        \REGS[18][21] ), .ZN(n1431) );
  OAI221_X1 U1035 ( .B1(n485), .B2(n143), .C1(n453), .C2(n139), .A(n1439), 
        .ZN(n1438) );
  AOI22_X1 U1036 ( .A1(n137), .A2(\REGS[3][21] ), .B1(n134), .B2(\REGS[2][21] ), .ZN(n1439) );
  OAI221_X1 U1037 ( .B1(n293), .B2(n2035), .C1(n290), .C2(n2003), .A(n777), 
        .ZN(n776) );
  AOI22_X1 U1038 ( .A1(\REGS[19][21] ), .A2(n287), .B1(\REGS[18][21] ), .B2(
        n284), .ZN(n777) );
  OAI221_X1 U1039 ( .B1(n245), .B2(n485), .C1(n242), .C2(n453), .A(n785), .ZN(
        n784) );
  AOI22_X1 U1040 ( .A1(\REGS[3][21] ), .A2(n239), .B1(\REGS[2][21] ), .B2(n236), .ZN(n785) );
  OAI221_X1 U1041 ( .B1(n2034), .B2(n191), .C1(n2002), .C2(n187), .A(n1449), 
        .ZN(n1448) );
  AOI22_X1 U1042 ( .A1(n185), .A2(\REGS[19][22] ), .B1(n182), .B2(
        \REGS[18][22] ), .ZN(n1449) );
  OAI221_X1 U1043 ( .B1(n484), .B2(n143), .C1(n452), .C2(n139), .A(n1457), 
        .ZN(n1456) );
  AOI22_X1 U1044 ( .A1(n137), .A2(\REGS[3][22] ), .B1(n134), .B2(\REGS[2][22] ), .ZN(n1457) );
  OAI221_X1 U1045 ( .B1(n293), .B2(n2034), .C1(n290), .C2(n2002), .A(n795), 
        .ZN(n794) );
  AOI22_X1 U1046 ( .A1(\REGS[19][22] ), .A2(n287), .B1(\REGS[18][22] ), .B2(
        n284), .ZN(n795) );
  OAI221_X1 U1047 ( .B1(n245), .B2(n484), .C1(n242), .C2(n452), .A(n803), .ZN(
        n802) );
  AOI22_X1 U1048 ( .A1(\REGS[3][22] ), .A2(n239), .B1(\REGS[2][22] ), .B2(n236), .ZN(n803) );
  OAI221_X1 U1049 ( .B1(n2033), .B2(n191), .C1(n2001), .C2(n187), .A(n1467), 
        .ZN(n1466) );
  AOI22_X1 U1050 ( .A1(n185), .A2(\REGS[19][23] ), .B1(n182), .B2(
        \REGS[18][23] ), .ZN(n1467) );
  OAI221_X1 U1051 ( .B1(n483), .B2(n143), .C1(n451), .C2(n139), .A(n1475), 
        .ZN(n1474) );
  AOI22_X1 U1052 ( .A1(n137), .A2(\REGS[3][23] ), .B1(n134), .B2(\REGS[2][23] ), .ZN(n1475) );
  OAI221_X1 U1053 ( .B1(n293), .B2(n2033), .C1(n290), .C2(n2001), .A(n813), 
        .ZN(n812) );
  AOI22_X1 U1054 ( .A1(\REGS[19][23] ), .A2(n287), .B1(\REGS[18][23] ), .B2(
        n284), .ZN(n813) );
  OAI221_X1 U1055 ( .B1(n245), .B2(n483), .C1(n242), .C2(n451), .A(n821), .ZN(
        n820) );
  AOI22_X1 U1056 ( .A1(\REGS[3][23] ), .A2(n239), .B1(\REGS[2][23] ), .B2(n236), .ZN(n821) );
  OAI221_X1 U1057 ( .B1(n2032), .B2(n191), .C1(n2000), .C2(n187), .A(n1485), 
        .ZN(n1484) );
  AOI22_X1 U1058 ( .A1(n185), .A2(\REGS[19][24] ), .B1(n182), .B2(
        \REGS[18][24] ), .ZN(n1485) );
  OAI221_X1 U1059 ( .B1(n482), .B2(n143), .C1(n450), .C2(n139), .A(n1493), 
        .ZN(n1492) );
  AOI22_X1 U1060 ( .A1(n137), .A2(\REGS[3][24] ), .B1(n134), .B2(\REGS[2][24] ), .ZN(n1493) );
  OAI221_X1 U1061 ( .B1(n293), .B2(n2032), .C1(n290), .C2(n2000), .A(n831), 
        .ZN(n830) );
  AOI22_X1 U1062 ( .A1(\REGS[19][24] ), .A2(n287), .B1(\REGS[18][24] ), .B2(
        n284), .ZN(n831) );
  OAI221_X1 U1063 ( .B1(n245), .B2(n482), .C1(n242), .C2(n450), .A(n839), .ZN(
        n838) );
  AOI22_X1 U1064 ( .A1(\REGS[3][24] ), .A2(n239), .B1(\REGS[2][24] ), .B2(n236), .ZN(n839) );
  OAI221_X1 U1065 ( .B1(n293), .B2(n2031), .C1(n290), .C2(n1999), .A(n849), 
        .ZN(n848) );
  AOI22_X1 U1066 ( .A1(\REGS[19][25] ), .A2(n287), .B1(\REGS[18][25] ), .B2(
        n284), .ZN(n849) );
  OAI221_X1 U1067 ( .B1(n245), .B2(n481), .C1(n242), .C2(n449), .A(n857), .ZN(
        n856) );
  AOI22_X1 U1068 ( .A1(\REGS[3][25] ), .A2(n239), .B1(\REGS[2][25] ), .B2(n236), .ZN(n857) );
  OAI221_X1 U1069 ( .B1(n293), .B2(n2030), .C1(n290), .C2(n1998), .A(n867), 
        .ZN(n866) );
  AOI22_X1 U1070 ( .A1(\REGS[19][26] ), .A2(n287), .B1(\REGS[18][26] ), .B2(
        n284), .ZN(n867) );
  OAI221_X1 U1071 ( .B1(n245), .B2(n480), .C1(n242), .C2(n448), .A(n875), .ZN(
        n874) );
  AOI22_X1 U1072 ( .A1(\REGS[3][26] ), .A2(n239), .B1(\REGS[2][26] ), .B2(n236), .ZN(n875) );
  OAI221_X1 U1073 ( .B1(n293), .B2(n2029), .C1(n290), .C2(n1997), .A(n885), 
        .ZN(n884) );
  AOI22_X1 U1074 ( .A1(\REGS[19][27] ), .A2(n287), .B1(\REGS[18][27] ), .B2(
        n284), .ZN(n885) );
  OAI221_X1 U1075 ( .B1(n245), .B2(n479), .C1(n242), .C2(n447), .A(n893), .ZN(
        n892) );
  AOI22_X1 U1076 ( .A1(\REGS[3][27] ), .A2(n239), .B1(\REGS[2][27] ), .B2(n236), .ZN(n893) );
  OAI221_X1 U1077 ( .B1(n293), .B2(n2028), .C1(n290), .C2(n1996), .A(n903), 
        .ZN(n902) );
  AOI22_X1 U1078 ( .A1(\REGS[19][28] ), .A2(n287), .B1(\REGS[18][28] ), .B2(
        n284), .ZN(n903) );
  OAI221_X1 U1079 ( .B1(n245), .B2(n478), .C1(n242), .C2(n446), .A(n911), .ZN(
        n910) );
  AOI22_X1 U1080 ( .A1(\REGS[3][28] ), .A2(n239), .B1(\REGS[2][28] ), .B2(n236), .ZN(n911) );
  OAI221_X1 U1081 ( .B1(n293), .B2(n2027), .C1(n290), .C2(n1995), .A(n921), 
        .ZN(n920) );
  AOI22_X1 U1082 ( .A1(\REGS[19][29] ), .A2(n287), .B1(\REGS[18][29] ), .B2(
        n284), .ZN(n921) );
  OAI221_X1 U1083 ( .B1(n245), .B2(n477), .C1(n242), .C2(n445), .A(n929), .ZN(
        n928) );
  AOI22_X1 U1084 ( .A1(\REGS[3][29] ), .A2(n239), .B1(\REGS[2][29] ), .B2(n236), .ZN(n929) );
  OAI221_X1 U1085 ( .B1(n293), .B2(n2026), .C1(n290), .C2(n1994), .A(n939), 
        .ZN(n938) );
  AOI22_X1 U1086 ( .A1(\REGS[19][30] ), .A2(n287), .B1(\REGS[18][30] ), .B2(
        n284), .ZN(n939) );
  OAI221_X1 U1087 ( .B1(n245), .B2(n476), .C1(n242), .C2(n444), .A(n947), .ZN(
        n946) );
  AOI22_X1 U1088 ( .A1(\REGS[3][30] ), .A2(n239), .B1(\REGS[2][30] ), .B2(n236), .ZN(n947) );
  OAI221_X1 U1089 ( .B1(n292), .B2(n2025), .C1(n289), .C2(n1993), .A(n957), 
        .ZN(n956) );
  AOI22_X1 U1090 ( .A1(\REGS[19][31] ), .A2(n286), .B1(\REGS[18][31] ), .B2(
        n283), .ZN(n957) );
  OAI221_X1 U1091 ( .B1(n244), .B2(n475), .C1(n241), .C2(n443), .A(n965), .ZN(
        n964) );
  AOI22_X1 U1092 ( .A1(\REGS[3][31] ), .A2(n238), .B1(\REGS[2][31] ), .B2(n235), .ZN(n965) );
  OAI221_X1 U1093 ( .B1(n282), .B2(n2109), .C1(n279), .C2(n2077), .A(n572), 
        .ZN(n563) );
  AOI22_X1 U1094 ( .A1(\REGS[23][11] ), .A2(n276), .B1(\REGS[22][11] ), .B2(
        n273), .ZN(n572) );
  OAI221_X1 U1095 ( .B1(n234), .B2(n1853), .C1(n231), .C2(n527), .A(n596), 
        .ZN(n587) );
  AOI22_X1 U1096 ( .A1(\REGS[7][11] ), .A2(n228), .B1(\REGS[6][11] ), .B2(n225), .ZN(n596) );
  OAI221_X1 U1097 ( .B1(n282), .B2(n2108), .C1(n279), .C2(n2076), .A(n616), 
        .ZN(n613) );
  AOI22_X1 U1098 ( .A1(\REGS[23][12] ), .A2(n276), .B1(\REGS[22][12] ), .B2(
        n273), .ZN(n616) );
  OAI221_X1 U1099 ( .B1(n234), .B2(n558), .C1(n231), .C2(n526), .A(n624), .ZN(
        n621) );
  AOI22_X1 U1100 ( .A1(\REGS[7][12] ), .A2(n228), .B1(\REGS[6][12] ), .B2(n225), .ZN(n624) );
  OAI221_X1 U1101 ( .B1(n282), .B2(n2107), .C1(n279), .C2(n2075), .A(n634), 
        .ZN(n631) );
  AOI22_X1 U1102 ( .A1(\REGS[23][13] ), .A2(n276), .B1(\REGS[22][13] ), .B2(
        n273), .ZN(n634) );
  OAI221_X1 U1103 ( .B1(n234), .B2(n557), .C1(n231), .C2(n525), .A(n642), .ZN(
        n639) );
  AOI22_X1 U1104 ( .A1(\REGS[7][13] ), .A2(n228), .B1(\REGS[6][13] ), .B2(n225), .ZN(n642) );
  OAI221_X1 U1105 ( .B1(n282), .B2(n2106), .C1(n279), .C2(n2074), .A(n652), 
        .ZN(n649) );
  AOI22_X1 U1106 ( .A1(\REGS[23][14] ), .A2(n276), .B1(\REGS[22][14] ), .B2(
        n273), .ZN(n652) );
  OAI221_X1 U1107 ( .B1(n234), .B2(n556), .C1(n231), .C2(n524), .A(n660), .ZN(
        n657) );
  AOI22_X1 U1108 ( .A1(\REGS[7][14] ), .A2(n228), .B1(\REGS[6][14] ), .B2(n225), .ZN(n660) );
  OAI221_X1 U1109 ( .B1(n282), .B2(n2105), .C1(n279), .C2(n2073), .A(n670), 
        .ZN(n667) );
  AOI22_X1 U1110 ( .A1(\REGS[23][15] ), .A2(n276), .B1(\REGS[22][15] ), .B2(
        n273), .ZN(n670) );
  OAI221_X1 U1111 ( .B1(n234), .B2(n555), .C1(n231), .C2(n523), .A(n678), .ZN(
        n675) );
  AOI22_X1 U1112 ( .A1(\REGS[7][15] ), .A2(n228), .B1(\REGS[6][15] ), .B2(n225), .ZN(n678) );
  OAI221_X1 U1113 ( .B1(n282), .B2(n2104), .C1(n279), .C2(n2072), .A(n688), 
        .ZN(n685) );
  AOI22_X1 U1114 ( .A1(\REGS[23][16] ), .A2(n276), .B1(\REGS[22][16] ), .B2(
        n273), .ZN(n688) );
  OAI221_X1 U1115 ( .B1(n234), .B2(n554), .C1(n231), .C2(n522), .A(n696), .ZN(
        n693) );
  AOI22_X1 U1116 ( .A1(\REGS[7][16] ), .A2(n228), .B1(\REGS[6][16] ), .B2(n225), .ZN(n696) );
  OAI221_X1 U1117 ( .B1(n282), .B2(n2103), .C1(n279), .C2(n2071), .A(n706), 
        .ZN(n703) );
  AOI22_X1 U1118 ( .A1(\REGS[23][17] ), .A2(n276), .B1(\REGS[22][17] ), .B2(
        n273), .ZN(n706) );
  OAI221_X1 U1119 ( .B1(n234), .B2(n553), .C1(n231), .C2(n521), .A(n714), .ZN(
        n711) );
  AOI22_X1 U1120 ( .A1(\REGS[7][17] ), .A2(n228), .B1(\REGS[6][17] ), .B2(n225), .ZN(n714) );
  OAI221_X1 U1121 ( .B1(n282), .B2(n2102), .C1(n279), .C2(n2070), .A(n724), 
        .ZN(n721) );
  AOI22_X1 U1122 ( .A1(\REGS[23][18] ), .A2(n276), .B1(\REGS[22][18] ), .B2(
        n273), .ZN(n724) );
  OAI221_X1 U1123 ( .B1(n234), .B2(n552), .C1(n231), .C2(n520), .A(n732), .ZN(
        n729) );
  AOI22_X1 U1124 ( .A1(\REGS[7][18] ), .A2(n228), .B1(\REGS[6][18] ), .B2(n225), .ZN(n732) );
  OAI221_X1 U1125 ( .B1(n2095), .B2(n180), .C1(n2063), .C2(n175), .A(n1504), 
        .ZN(n1501) );
  AOI22_X1 U1126 ( .A1(n174), .A2(\REGS[23][25] ), .B1(n171), .B2(
        \REGS[22][25] ), .ZN(n1504) );
  OAI221_X1 U1127 ( .B1(n545), .B2(n132), .C1(n513), .C2(n127), .A(n1512), 
        .ZN(n1509) );
  AOI22_X1 U1128 ( .A1(n126), .A2(\REGS[7][25] ), .B1(n123), .B2(\REGS[6][25] ), .ZN(n1512) );
  OAI221_X1 U1129 ( .B1(n2094), .B2(n180), .C1(n2062), .C2(n175), .A(n1522), 
        .ZN(n1519) );
  AOI22_X1 U1130 ( .A1(n174), .A2(\REGS[23][26] ), .B1(n171), .B2(
        \REGS[22][26] ), .ZN(n1522) );
  OAI221_X1 U1131 ( .B1(n544), .B2(n132), .C1(n512), .C2(n127), .A(n1530), 
        .ZN(n1527) );
  AOI22_X1 U1132 ( .A1(n126), .A2(\REGS[7][26] ), .B1(n123), .B2(\REGS[6][26] ), .ZN(n1530) );
  OAI221_X1 U1133 ( .B1(n2093), .B2(n180), .C1(n2061), .C2(n175), .A(n1540), 
        .ZN(n1537) );
  AOI22_X1 U1134 ( .A1(n174), .A2(\REGS[23][27] ), .B1(n171), .B2(
        \REGS[22][27] ), .ZN(n1540) );
  OAI221_X1 U1135 ( .B1(n543), .B2(n132), .C1(n511), .C2(n127), .A(n1548), 
        .ZN(n1545) );
  AOI22_X1 U1136 ( .A1(n126), .A2(\REGS[7][27] ), .B1(n123), .B2(\REGS[6][27] ), .ZN(n1548) );
  OAI221_X1 U1137 ( .B1(n2092), .B2(n180), .C1(n2060), .C2(n175), .A(n1558), 
        .ZN(n1555) );
  AOI22_X1 U1138 ( .A1(n174), .A2(\REGS[23][28] ), .B1(n171), .B2(
        \REGS[22][28] ), .ZN(n1558) );
  OAI221_X1 U1139 ( .B1(n542), .B2(n132), .C1(n510), .C2(n127), .A(n1566), 
        .ZN(n1563) );
  AOI22_X1 U1140 ( .A1(n126), .A2(\REGS[7][28] ), .B1(n123), .B2(\REGS[6][28] ), .ZN(n1566) );
  OAI221_X1 U1141 ( .B1(n2091), .B2(n180), .C1(n2059), .C2(n175), .A(n1576), 
        .ZN(n1573) );
  AOI22_X1 U1142 ( .A1(n174), .A2(\REGS[23][29] ), .B1(n171), .B2(
        \REGS[22][29] ), .ZN(n1576) );
  OAI221_X1 U1143 ( .B1(n541), .B2(n132), .C1(n509), .C2(n127), .A(n1584), 
        .ZN(n1581) );
  AOI22_X1 U1144 ( .A1(n126), .A2(\REGS[7][29] ), .B1(n123), .B2(\REGS[6][29] ), .ZN(n1584) );
  OAI221_X1 U1145 ( .B1(n2090), .B2(n180), .C1(n2058), .C2(n175), .A(n1594), 
        .ZN(n1591) );
  AOI22_X1 U1146 ( .A1(n174), .A2(\REGS[23][30] ), .B1(n171), .B2(
        \REGS[22][30] ), .ZN(n1594) );
  OAI221_X1 U1147 ( .B1(n540), .B2(n132), .C1(n508), .C2(n127), .A(n1602), 
        .ZN(n1599) );
  AOI22_X1 U1148 ( .A1(n126), .A2(\REGS[7][30] ), .B1(n123), .B2(\REGS[6][30] ), .ZN(n1602) );
  OAI221_X1 U1149 ( .B1(n2089), .B2(n180), .C1(n2057), .C2(n175), .A(n1616), 
        .ZN(n1609) );
  AOI22_X1 U1150 ( .A1(n174), .A2(\REGS[23][31] ), .B1(n171), .B2(
        \REGS[22][31] ), .ZN(n1616) );
  OAI221_X1 U1151 ( .B1(n539), .B2(n132), .C1(n507), .C2(n127), .A(n1632), 
        .ZN(n1627) );
  AOI22_X1 U1152 ( .A1(n126), .A2(\REGS[7][31] ), .B1(n123), .B2(\REGS[6][31] ), .ZN(n1632) );
  OAI221_X1 U1153 ( .B1(n280), .B2(n2120), .C1(n277), .C2(n2088), .A(n1646), 
        .ZN(n1643) );
  AOI22_X1 U1154 ( .A1(\REGS[23][0] ), .A2(n274), .B1(\REGS[22][0] ), .B2(n271), .ZN(n1646) );
  OAI221_X1 U1155 ( .B1(n232), .B2(n1864), .C1(n229), .C2(n538), .A(n1654), 
        .ZN(n1651) );
  AOI22_X1 U1156 ( .A1(\REGS[7][0] ), .A2(n226), .B1(\REGS[6][0] ), .B2(n223), 
        .ZN(n1654) );
  OAI221_X1 U1157 ( .B1(n178), .B2(n2120), .C1(n177), .C2(n2088), .A(n1028), 
        .ZN(n1019) );
  AOI22_X1 U1158 ( .A1(\REGS[23][0] ), .A2(n172), .B1(\REGS[22][0] ), .B2(n169), .ZN(n1028) );
  OAI221_X1 U1159 ( .B1(n130), .B2(n1864), .C1(n129), .C2(n538), .A(n1052), 
        .ZN(n1043) );
  AOI22_X1 U1160 ( .A1(\REGS[7][0] ), .A2(n124), .B1(\REGS[6][0] ), .B2(n121), 
        .ZN(n1052) );
  OAI221_X1 U1161 ( .B1(n280), .B2(n2119), .C1(n277), .C2(n2087), .A(n1664), 
        .ZN(n1661) );
  AOI22_X1 U1162 ( .A1(\REGS[23][1] ), .A2(n274), .B1(\REGS[22][1] ), .B2(n271), .ZN(n1664) );
  OAI221_X1 U1163 ( .B1(n232), .B2(n1863), .C1(n229), .C2(n537), .A(n1672), 
        .ZN(n1669) );
  AOI22_X1 U1164 ( .A1(\REGS[7][1] ), .A2(n226), .B1(\REGS[6][1] ), .B2(n223), 
        .ZN(n1672) );
  OAI221_X1 U1165 ( .B1(n178), .B2(n2119), .C1(n177), .C2(n2087), .A(n1072), 
        .ZN(n1069) );
  AOI22_X1 U1166 ( .A1(\REGS[23][1] ), .A2(n172), .B1(\REGS[22][1] ), .B2(n169), .ZN(n1072) );
  OAI221_X1 U1167 ( .B1(n130), .B2(n1863), .C1(n129), .C2(n537), .A(n1080), 
        .ZN(n1077) );
  AOI22_X1 U1168 ( .A1(\REGS[7][1] ), .A2(n124), .B1(\REGS[6][1] ), .B2(n121), 
        .ZN(n1080) );
  OAI221_X1 U1169 ( .B1(n280), .B2(n2118), .C1(n277), .C2(n2086), .A(n1682), 
        .ZN(n1679) );
  AOI22_X1 U1170 ( .A1(\REGS[23][2] ), .A2(n274), .B1(\REGS[22][2] ), .B2(n271), .ZN(n1682) );
  OAI221_X1 U1171 ( .B1(n232), .B2(n1862), .C1(n229), .C2(n536), .A(n1690), 
        .ZN(n1687) );
  AOI22_X1 U1172 ( .A1(\REGS[7][2] ), .A2(n226), .B1(\REGS[6][2] ), .B2(n223), 
        .ZN(n1690) );
  OAI221_X1 U1173 ( .B1(n178), .B2(n2118), .C1(n177), .C2(n2086), .A(n1090), 
        .ZN(n1087) );
  AOI22_X1 U1174 ( .A1(\REGS[23][2] ), .A2(n172), .B1(\REGS[22][2] ), .B2(n169), .ZN(n1090) );
  OAI221_X1 U1175 ( .B1(n130), .B2(n1862), .C1(n129), .C2(n536), .A(n1098), 
        .ZN(n1095) );
  AOI22_X1 U1176 ( .A1(\REGS[7][2] ), .A2(n124), .B1(\REGS[6][2] ), .B2(n121), 
        .ZN(n1098) );
  OAI221_X1 U1177 ( .B1(n280), .B2(n2117), .C1(n277), .C2(n2085), .A(n1700), 
        .ZN(n1697) );
  AOI22_X1 U1178 ( .A1(\REGS[23][3] ), .A2(n274), .B1(\REGS[22][3] ), .B2(n271), .ZN(n1700) );
  OAI221_X1 U1179 ( .B1(n232), .B2(n1861), .C1(n229), .C2(n535), .A(n1708), 
        .ZN(n1705) );
  AOI22_X1 U1180 ( .A1(\REGS[7][3] ), .A2(n226), .B1(\REGS[6][3] ), .B2(n223), 
        .ZN(n1708) );
  OAI221_X1 U1181 ( .B1(n178), .B2(n2117), .C1(n177), .C2(n2085), .A(n1108), 
        .ZN(n1105) );
  AOI22_X1 U1182 ( .A1(\REGS[23][3] ), .A2(n172), .B1(\REGS[22][3] ), .B2(n169), .ZN(n1108) );
  OAI221_X1 U1183 ( .B1(n130), .B2(n1861), .C1(n129), .C2(n535), .A(n1116), 
        .ZN(n1113) );
  AOI22_X1 U1184 ( .A1(\REGS[7][3] ), .A2(n124), .B1(\REGS[6][3] ), .B2(n121), 
        .ZN(n1116) );
  OAI221_X1 U1185 ( .B1(n280), .B2(n2116), .C1(n277), .C2(n2084), .A(n1718), 
        .ZN(n1715) );
  AOI22_X1 U1186 ( .A1(\REGS[23][4] ), .A2(n274), .B1(\REGS[22][4] ), .B2(n271), .ZN(n1718) );
  OAI221_X1 U1187 ( .B1(n232), .B2(n1860), .C1(n229), .C2(n534), .A(n1726), 
        .ZN(n1723) );
  AOI22_X1 U1188 ( .A1(\REGS[7][4] ), .A2(n226), .B1(\REGS[6][4] ), .B2(n223), 
        .ZN(n1726) );
  OAI221_X1 U1189 ( .B1(n178), .B2(n2116), .C1(n177), .C2(n2084), .A(n1126), 
        .ZN(n1123) );
  AOI22_X1 U1190 ( .A1(\REGS[23][4] ), .A2(n172), .B1(\REGS[22][4] ), .B2(n169), .ZN(n1126) );
  OAI221_X1 U1191 ( .B1(n130), .B2(n1860), .C1(n129), .C2(n534), .A(n1134), 
        .ZN(n1131) );
  AOI22_X1 U1192 ( .A1(\REGS[7][4] ), .A2(n124), .B1(\REGS[6][4] ), .B2(n121), 
        .ZN(n1134) );
  OAI221_X1 U1193 ( .B1(n280), .B2(n2115), .C1(n277), .C2(n2083), .A(n1736), 
        .ZN(n1733) );
  AOI22_X1 U1194 ( .A1(\REGS[23][5] ), .A2(n274), .B1(\REGS[22][5] ), .B2(n271), .ZN(n1736) );
  OAI221_X1 U1195 ( .B1(n232), .B2(n1859), .C1(n229), .C2(n533), .A(n1744), 
        .ZN(n1741) );
  AOI22_X1 U1196 ( .A1(\REGS[7][5] ), .A2(n226), .B1(\REGS[6][5] ), .B2(n223), 
        .ZN(n1744) );
  OAI221_X1 U1197 ( .B1(n178), .B2(n2115), .C1(n177), .C2(n2083), .A(n1144), 
        .ZN(n1141) );
  AOI22_X1 U1198 ( .A1(\REGS[23][5] ), .A2(n172), .B1(\REGS[22][5] ), .B2(n169), .ZN(n1144) );
  OAI221_X1 U1199 ( .B1(n130), .B2(n1859), .C1(n129), .C2(n533), .A(n1152), 
        .ZN(n1149) );
  AOI22_X1 U1200 ( .A1(\REGS[7][5] ), .A2(n124), .B1(\REGS[6][5] ), .B2(n121), 
        .ZN(n1152) );
  OAI221_X1 U1201 ( .B1(n280), .B2(n2114), .C1(n277), .C2(n2082), .A(n1754), 
        .ZN(n1751) );
  AOI22_X1 U1202 ( .A1(\REGS[23][6] ), .A2(n274), .B1(\REGS[22][6] ), .B2(n271), .ZN(n1754) );
  OAI221_X1 U1203 ( .B1(n232), .B2(n1858), .C1(n229), .C2(n532), .A(n1762), 
        .ZN(n1759) );
  AOI22_X1 U1204 ( .A1(\REGS[7][6] ), .A2(n226), .B1(\REGS[6][6] ), .B2(n223), 
        .ZN(n1762) );
  OAI221_X1 U1205 ( .B1(n178), .B2(n2114), .C1(n177), .C2(n2082), .A(n1162), 
        .ZN(n1159) );
  AOI22_X1 U1206 ( .A1(\REGS[23][6] ), .A2(n172), .B1(\REGS[22][6] ), .B2(n169), .ZN(n1162) );
  OAI221_X1 U1207 ( .B1(n130), .B2(n1858), .C1(n129), .C2(n532), .A(n1170), 
        .ZN(n1167) );
  AOI22_X1 U1208 ( .A1(\REGS[7][6] ), .A2(n124), .B1(\REGS[6][6] ), .B2(n121), 
        .ZN(n1170) );
  OAI221_X1 U1209 ( .B1(n280), .B2(n2113), .C1(n277), .C2(n2081), .A(n1772), 
        .ZN(n1769) );
  AOI22_X1 U1210 ( .A1(\REGS[23][7] ), .A2(n274), .B1(\REGS[22][7] ), .B2(n271), .ZN(n1772) );
  OAI221_X1 U1211 ( .B1(n232), .B2(n1857), .C1(n229), .C2(n531), .A(n1780), 
        .ZN(n1777) );
  AOI22_X1 U1212 ( .A1(\REGS[7][7] ), .A2(n226), .B1(\REGS[6][7] ), .B2(n223), 
        .ZN(n1780) );
  OAI221_X1 U1213 ( .B1(n178), .B2(n2113), .C1(n177), .C2(n2081), .A(n1180), 
        .ZN(n1177) );
  AOI22_X1 U1214 ( .A1(\REGS[23][7] ), .A2(n172), .B1(\REGS[22][7] ), .B2(n169), .ZN(n1180) );
  OAI221_X1 U1215 ( .B1(n130), .B2(n1857), .C1(n129), .C2(n531), .A(n1188), 
        .ZN(n1185) );
  AOI22_X1 U1216 ( .A1(\REGS[7][7] ), .A2(n124), .B1(\REGS[6][7] ), .B2(n121), 
        .ZN(n1188) );
  OAI221_X1 U1217 ( .B1(n280), .B2(n2112), .C1(n277), .C2(n2080), .A(n1790), 
        .ZN(n1787) );
  AOI22_X1 U1218 ( .A1(\REGS[23][8] ), .A2(n274), .B1(\REGS[22][8] ), .B2(n271), .ZN(n1790) );
  OAI221_X1 U1219 ( .B1(n232), .B2(n1856), .C1(n229), .C2(n530), .A(n1798), 
        .ZN(n1795) );
  AOI22_X1 U1220 ( .A1(\REGS[7][8] ), .A2(n226), .B1(\REGS[6][8] ), .B2(n223), 
        .ZN(n1798) );
  OAI221_X1 U1221 ( .B1(n178), .B2(n2112), .C1(n176), .C2(n2080), .A(n1198), 
        .ZN(n1195) );
  AOI22_X1 U1222 ( .A1(\REGS[23][8] ), .A2(n172), .B1(\REGS[22][8] ), .B2(n169), .ZN(n1198) );
  OAI221_X1 U1223 ( .B1(n130), .B2(n1856), .C1(n128), .C2(n530), .A(n1206), 
        .ZN(n1203) );
  AOI22_X1 U1224 ( .A1(\REGS[7][8] ), .A2(n124), .B1(\REGS[6][8] ), .B2(n121), 
        .ZN(n1206) );
  OAI221_X1 U1225 ( .B1(n280), .B2(n2111), .C1(n277), .C2(n2079), .A(n1808), 
        .ZN(n1805) );
  AOI22_X1 U1226 ( .A1(\REGS[23][9] ), .A2(n274), .B1(\REGS[22][9] ), .B2(n271), .ZN(n1808) );
  OAI221_X1 U1227 ( .B1(n232), .B2(n1855), .C1(n229), .C2(n529), .A(n1816), 
        .ZN(n1813) );
  AOI22_X1 U1228 ( .A1(\REGS[7][9] ), .A2(n226), .B1(\REGS[6][9] ), .B2(n223), 
        .ZN(n1816) );
  OAI221_X1 U1229 ( .B1(n178), .B2(n2111), .C1(n176), .C2(n2079), .A(n1216), 
        .ZN(n1213) );
  AOI22_X1 U1230 ( .A1(\REGS[23][9] ), .A2(n172), .B1(\REGS[22][9] ), .B2(n169), .ZN(n1216) );
  OAI221_X1 U1231 ( .B1(n130), .B2(n1855), .C1(n128), .C2(n529), .A(n1224), 
        .ZN(n1221) );
  AOI22_X1 U1232 ( .A1(\REGS[7][9] ), .A2(n124), .B1(\REGS[6][9] ), .B2(n121), 
        .ZN(n1224) );
  OAI221_X1 U1233 ( .B1(n280), .B2(n2110), .C1(n277), .C2(n2078), .A(n1830), 
        .ZN(n1823) );
  AOI22_X1 U1234 ( .A1(\REGS[23][10] ), .A2(n274), .B1(\REGS[22][10] ), .B2(
        n271), .ZN(n1830) );
  OAI221_X1 U1235 ( .B1(n232), .B2(n1854), .C1(n229), .C2(n528), .A(n1846), 
        .ZN(n1841) );
  AOI22_X1 U1236 ( .A1(\REGS[7][10] ), .A2(n226), .B1(\REGS[6][10] ), .B2(n223), .ZN(n1846) );
  OAI221_X1 U1237 ( .B1(n178), .B2(n2110), .C1(n176), .C2(n2078), .A(n1234), 
        .ZN(n1231) );
  AOI22_X1 U1238 ( .A1(\REGS[23][10] ), .A2(n172), .B1(\REGS[22][10] ), .B2(
        n169), .ZN(n1234) );
  OAI221_X1 U1239 ( .B1(n130), .B2(n1854), .C1(n128), .C2(n528), .A(n1242), 
        .ZN(n1239) );
  AOI22_X1 U1240 ( .A1(\REGS[7][10] ), .A2(n124), .B1(\REGS[6][10] ), .B2(n121), .ZN(n1242) );
  OAI221_X1 U1241 ( .B1(n2109), .B2(n178), .C1(n2077), .C2(n176), .A(n1252), 
        .ZN(n1249) );
  AOI22_X1 U1242 ( .A1(n172), .A2(\REGS[23][11] ), .B1(n169), .B2(
        \REGS[22][11] ), .ZN(n1252) );
  OAI221_X1 U1243 ( .B1(n1853), .B2(n130), .C1(n527), .C2(n128), .A(n1260), 
        .ZN(n1257) );
  AOI22_X1 U1244 ( .A1(n124), .A2(\REGS[7][11] ), .B1(n121), .B2(\REGS[6][11] ), .ZN(n1260) );
  OAI221_X1 U1245 ( .B1(n2108), .B2(n179), .C1(n2076), .C2(n176), .A(n1270), 
        .ZN(n1267) );
  AOI22_X1 U1246 ( .A1(n173), .A2(\REGS[23][12] ), .B1(n170), .B2(
        \REGS[22][12] ), .ZN(n1270) );
  OAI221_X1 U1247 ( .B1(n558), .B2(n131), .C1(n526), .C2(n128), .A(n1278), 
        .ZN(n1275) );
  AOI22_X1 U1248 ( .A1(n125), .A2(\REGS[7][12] ), .B1(n122), .B2(\REGS[6][12] ), .ZN(n1278) );
  OAI221_X1 U1249 ( .B1(n2107), .B2(n179), .C1(n2075), .C2(n176), .A(n1288), 
        .ZN(n1285) );
  AOI22_X1 U1250 ( .A1(n173), .A2(\REGS[23][13] ), .B1(n170), .B2(
        \REGS[22][13] ), .ZN(n1288) );
  OAI221_X1 U1251 ( .B1(n557), .B2(n131), .C1(n525), .C2(n128), .A(n1296), 
        .ZN(n1293) );
  AOI22_X1 U1252 ( .A1(n125), .A2(\REGS[7][13] ), .B1(n122), .B2(\REGS[6][13] ), .ZN(n1296) );
  OAI221_X1 U1253 ( .B1(n2106), .B2(n179), .C1(n2074), .C2(n176), .A(n1306), 
        .ZN(n1303) );
  AOI22_X1 U1254 ( .A1(n173), .A2(\REGS[23][14] ), .B1(n170), .B2(
        \REGS[22][14] ), .ZN(n1306) );
  OAI221_X1 U1255 ( .B1(n556), .B2(n131), .C1(n524), .C2(n128), .A(n1314), 
        .ZN(n1311) );
  AOI22_X1 U1256 ( .A1(n125), .A2(\REGS[7][14] ), .B1(n122), .B2(\REGS[6][14] ), .ZN(n1314) );
  OAI221_X1 U1257 ( .B1(n2105), .B2(n179), .C1(n2073), .C2(n176), .A(n1324), 
        .ZN(n1321) );
  AOI22_X1 U1258 ( .A1(n173), .A2(\REGS[23][15] ), .B1(n170), .B2(
        \REGS[22][15] ), .ZN(n1324) );
  OAI221_X1 U1259 ( .B1(n555), .B2(n131), .C1(n523), .C2(n128), .A(n1332), 
        .ZN(n1329) );
  AOI22_X1 U1260 ( .A1(n125), .A2(\REGS[7][15] ), .B1(n122), .B2(\REGS[6][15] ), .ZN(n1332) );
  OAI221_X1 U1261 ( .B1(n2104), .B2(n179), .C1(n2072), .C2(n176), .A(n1342), 
        .ZN(n1339) );
  AOI22_X1 U1262 ( .A1(n173), .A2(\REGS[23][16] ), .B1(n170), .B2(
        \REGS[22][16] ), .ZN(n1342) );
  OAI221_X1 U1263 ( .B1(n554), .B2(n131), .C1(n522), .C2(n128), .A(n1350), 
        .ZN(n1347) );
  AOI22_X1 U1264 ( .A1(n125), .A2(\REGS[7][16] ), .B1(n122), .B2(\REGS[6][16] ), .ZN(n1350) );
  OAI221_X1 U1265 ( .B1(n2103), .B2(n179), .C1(n2071), .C2(n176), .A(n1360), 
        .ZN(n1357) );
  AOI22_X1 U1266 ( .A1(n173), .A2(\REGS[23][17] ), .B1(n170), .B2(
        \REGS[22][17] ), .ZN(n1360) );
  OAI221_X1 U1267 ( .B1(n553), .B2(n131), .C1(n521), .C2(n128), .A(n1368), 
        .ZN(n1365) );
  AOI22_X1 U1268 ( .A1(n125), .A2(\REGS[7][17] ), .B1(n122), .B2(\REGS[6][17] ), .ZN(n1368) );
  OAI221_X1 U1269 ( .B1(n2102), .B2(n179), .C1(n2070), .C2(n176), .A(n1378), 
        .ZN(n1375) );
  AOI22_X1 U1270 ( .A1(n173), .A2(\REGS[23][18] ), .B1(n170), .B2(
        \REGS[22][18] ), .ZN(n1378) );
  OAI221_X1 U1271 ( .B1(n552), .B2(n131), .C1(n520), .C2(n128), .A(n1386), 
        .ZN(n1383) );
  AOI22_X1 U1272 ( .A1(n125), .A2(\REGS[7][18] ), .B1(n122), .B2(\REGS[6][18] ), .ZN(n1386) );
  OAI221_X1 U1273 ( .B1(n2101), .B2(n179), .C1(n2069), .C2(n176), .A(n1396), 
        .ZN(n1393) );
  AOI22_X1 U1274 ( .A1(n173), .A2(\REGS[23][19] ), .B1(n170), .B2(
        \REGS[22][19] ), .ZN(n1396) );
  OAI221_X1 U1275 ( .B1(n551), .B2(n131), .C1(n519), .C2(n128), .A(n1404), 
        .ZN(n1401) );
  AOI22_X1 U1276 ( .A1(n125), .A2(\REGS[7][19] ), .B1(n122), .B2(\REGS[6][19] ), .ZN(n1404) );
  OAI221_X1 U1277 ( .B1(n281), .B2(n2101), .C1(n278), .C2(n2069), .A(n742), 
        .ZN(n739) );
  AOI22_X1 U1278 ( .A1(\REGS[23][19] ), .A2(n275), .B1(\REGS[22][19] ), .B2(
        n272), .ZN(n742) );
  OAI221_X1 U1279 ( .B1(n233), .B2(n551), .C1(n230), .C2(n519), .A(n750), .ZN(
        n747) );
  AOI22_X1 U1280 ( .A1(\REGS[7][19] ), .A2(n227), .B1(\REGS[6][19] ), .B2(n224), .ZN(n750) );
  OAI221_X1 U1281 ( .B1(n2100), .B2(n179), .C1(n2068), .C2(n175), .A(n1414), 
        .ZN(n1411) );
  AOI22_X1 U1282 ( .A1(n173), .A2(\REGS[23][20] ), .B1(n170), .B2(
        \REGS[22][20] ), .ZN(n1414) );
  OAI221_X1 U1283 ( .B1(n550), .B2(n131), .C1(n518), .C2(n127), .A(n1422), 
        .ZN(n1419) );
  AOI22_X1 U1284 ( .A1(n125), .A2(\REGS[7][20] ), .B1(n122), .B2(\REGS[6][20] ), .ZN(n1422) );
  OAI221_X1 U1285 ( .B1(n281), .B2(n2100), .C1(n278), .C2(n2068), .A(n760), 
        .ZN(n757) );
  AOI22_X1 U1286 ( .A1(\REGS[23][20] ), .A2(n275), .B1(\REGS[22][20] ), .B2(
        n272), .ZN(n760) );
  OAI221_X1 U1287 ( .B1(n233), .B2(n550), .C1(n230), .C2(n518), .A(n768), .ZN(
        n765) );
  AOI22_X1 U1288 ( .A1(\REGS[7][20] ), .A2(n227), .B1(\REGS[6][20] ), .B2(n224), .ZN(n768) );
  OAI221_X1 U1289 ( .B1(n2099), .B2(n179), .C1(n2067), .C2(n175), .A(n1432), 
        .ZN(n1429) );
  AOI22_X1 U1290 ( .A1(n173), .A2(\REGS[23][21] ), .B1(n170), .B2(
        \REGS[22][21] ), .ZN(n1432) );
  OAI221_X1 U1291 ( .B1(n549), .B2(n131), .C1(n517), .C2(n127), .A(n1440), 
        .ZN(n1437) );
  AOI22_X1 U1292 ( .A1(n125), .A2(\REGS[7][21] ), .B1(n122), .B2(\REGS[6][21] ), .ZN(n1440) );
  OAI221_X1 U1293 ( .B1(n281), .B2(n2099), .C1(n278), .C2(n2067), .A(n778), 
        .ZN(n775) );
  AOI22_X1 U1294 ( .A1(\REGS[23][21] ), .A2(n275), .B1(\REGS[22][21] ), .B2(
        n272), .ZN(n778) );
  OAI221_X1 U1295 ( .B1(n233), .B2(n549), .C1(n230), .C2(n517), .A(n786), .ZN(
        n783) );
  AOI22_X1 U1296 ( .A1(\REGS[7][21] ), .A2(n227), .B1(\REGS[6][21] ), .B2(n224), .ZN(n786) );
  OAI221_X1 U1297 ( .B1(n2098), .B2(n179), .C1(n2066), .C2(n175), .A(n1450), 
        .ZN(n1447) );
  AOI22_X1 U1298 ( .A1(n173), .A2(\REGS[23][22] ), .B1(n170), .B2(
        \REGS[22][22] ), .ZN(n1450) );
  OAI221_X1 U1299 ( .B1(n548), .B2(n131), .C1(n516), .C2(n127), .A(n1458), 
        .ZN(n1455) );
  AOI22_X1 U1300 ( .A1(n125), .A2(\REGS[7][22] ), .B1(n122), .B2(\REGS[6][22] ), .ZN(n1458) );
  OAI221_X1 U1301 ( .B1(n281), .B2(n2098), .C1(n278), .C2(n2066), .A(n796), 
        .ZN(n793) );
  AOI22_X1 U1302 ( .A1(\REGS[23][22] ), .A2(n275), .B1(\REGS[22][22] ), .B2(
        n272), .ZN(n796) );
  OAI221_X1 U1303 ( .B1(n233), .B2(n548), .C1(n230), .C2(n516), .A(n804), .ZN(
        n801) );
  AOI22_X1 U1304 ( .A1(\REGS[7][22] ), .A2(n227), .B1(\REGS[6][22] ), .B2(n224), .ZN(n804) );
  OAI221_X1 U1305 ( .B1(n2097), .B2(n179), .C1(n2065), .C2(n175), .A(n1468), 
        .ZN(n1465) );
  AOI22_X1 U1306 ( .A1(n173), .A2(\REGS[23][23] ), .B1(n170), .B2(
        \REGS[22][23] ), .ZN(n1468) );
  OAI221_X1 U1307 ( .B1(n547), .B2(n131), .C1(n515), .C2(n127), .A(n1476), 
        .ZN(n1473) );
  AOI22_X1 U1308 ( .A1(n125), .A2(\REGS[7][23] ), .B1(n122), .B2(\REGS[6][23] ), .ZN(n1476) );
  OAI221_X1 U1309 ( .B1(n281), .B2(n2097), .C1(n278), .C2(n2065), .A(n814), 
        .ZN(n811) );
  AOI22_X1 U1310 ( .A1(\REGS[23][23] ), .A2(n275), .B1(\REGS[22][23] ), .B2(
        n272), .ZN(n814) );
  OAI221_X1 U1311 ( .B1(n233), .B2(n547), .C1(n230), .C2(n515), .A(n822), .ZN(
        n819) );
  AOI22_X1 U1312 ( .A1(\REGS[7][23] ), .A2(n227), .B1(\REGS[6][23] ), .B2(n224), .ZN(n822) );
  OAI221_X1 U1313 ( .B1(n2096), .B2(n179), .C1(n2064), .C2(n175), .A(n1486), 
        .ZN(n1483) );
  AOI22_X1 U1314 ( .A1(n173), .A2(\REGS[23][24] ), .B1(n170), .B2(
        \REGS[22][24] ), .ZN(n1486) );
  OAI221_X1 U1315 ( .B1(n546), .B2(n131), .C1(n514), .C2(n127), .A(n1494), 
        .ZN(n1491) );
  AOI22_X1 U1316 ( .A1(n125), .A2(\REGS[7][24] ), .B1(n122), .B2(\REGS[6][24] ), .ZN(n1494) );
  OAI221_X1 U1317 ( .B1(n281), .B2(n2096), .C1(n278), .C2(n2064), .A(n832), 
        .ZN(n829) );
  AOI22_X1 U1318 ( .A1(\REGS[23][24] ), .A2(n275), .B1(\REGS[22][24] ), .B2(
        n272), .ZN(n832) );
  OAI221_X1 U1319 ( .B1(n233), .B2(n546), .C1(n230), .C2(n514), .A(n840), .ZN(
        n837) );
  AOI22_X1 U1320 ( .A1(\REGS[7][24] ), .A2(n227), .B1(\REGS[6][24] ), .B2(n224), .ZN(n840) );
  OAI221_X1 U1321 ( .B1(n281), .B2(n2095), .C1(n278), .C2(n2063), .A(n850), 
        .ZN(n847) );
  AOI22_X1 U1322 ( .A1(\REGS[23][25] ), .A2(n275), .B1(\REGS[22][25] ), .B2(
        n272), .ZN(n850) );
  OAI221_X1 U1323 ( .B1(n233), .B2(n545), .C1(n230), .C2(n513), .A(n858), .ZN(
        n855) );
  AOI22_X1 U1324 ( .A1(\REGS[7][25] ), .A2(n227), .B1(\REGS[6][25] ), .B2(n224), .ZN(n858) );
  OAI221_X1 U1325 ( .B1(n281), .B2(n2094), .C1(n278), .C2(n2062), .A(n868), 
        .ZN(n865) );
  AOI22_X1 U1326 ( .A1(\REGS[23][26] ), .A2(n275), .B1(\REGS[22][26] ), .B2(
        n272), .ZN(n868) );
  OAI221_X1 U1327 ( .B1(n233), .B2(n544), .C1(n230), .C2(n512), .A(n876), .ZN(
        n873) );
  AOI22_X1 U1328 ( .A1(\REGS[7][26] ), .A2(n227), .B1(\REGS[6][26] ), .B2(n224), .ZN(n876) );
  OAI221_X1 U1329 ( .B1(n281), .B2(n2093), .C1(n278), .C2(n2061), .A(n886), 
        .ZN(n883) );
  AOI22_X1 U1330 ( .A1(\REGS[23][27] ), .A2(n275), .B1(\REGS[22][27] ), .B2(
        n272), .ZN(n886) );
  OAI221_X1 U1331 ( .B1(n233), .B2(n543), .C1(n230), .C2(n511), .A(n894), .ZN(
        n891) );
  AOI22_X1 U1332 ( .A1(\REGS[7][27] ), .A2(n227), .B1(\REGS[6][27] ), .B2(n224), .ZN(n894) );
  OAI221_X1 U1333 ( .B1(n281), .B2(n2092), .C1(n278), .C2(n2060), .A(n904), 
        .ZN(n901) );
  AOI22_X1 U1334 ( .A1(\REGS[23][28] ), .A2(n275), .B1(\REGS[22][28] ), .B2(
        n272), .ZN(n904) );
  OAI221_X1 U1335 ( .B1(n233), .B2(n542), .C1(n230), .C2(n510), .A(n912), .ZN(
        n909) );
  AOI22_X1 U1336 ( .A1(\REGS[7][28] ), .A2(n227), .B1(\REGS[6][28] ), .B2(n224), .ZN(n912) );
  OAI221_X1 U1337 ( .B1(n281), .B2(n2091), .C1(n278), .C2(n2059), .A(n922), 
        .ZN(n919) );
  AOI22_X1 U1338 ( .A1(\REGS[23][29] ), .A2(n275), .B1(\REGS[22][29] ), .B2(
        n272), .ZN(n922) );
  OAI221_X1 U1339 ( .B1(n233), .B2(n541), .C1(n230), .C2(n509), .A(n930), .ZN(
        n927) );
  AOI22_X1 U1340 ( .A1(\REGS[7][29] ), .A2(n227), .B1(\REGS[6][29] ), .B2(n224), .ZN(n930) );
  OAI221_X1 U1341 ( .B1(n281), .B2(n2090), .C1(n278), .C2(n2058), .A(n940), 
        .ZN(n937) );
  AOI22_X1 U1342 ( .A1(\REGS[23][30] ), .A2(n275), .B1(\REGS[22][30] ), .B2(
        n272), .ZN(n940) );
  OAI221_X1 U1343 ( .B1(n233), .B2(n540), .C1(n230), .C2(n508), .A(n948), .ZN(
        n945) );
  AOI22_X1 U1344 ( .A1(\REGS[7][30] ), .A2(n227), .B1(\REGS[6][30] ), .B2(n224), .ZN(n948) );
  OAI221_X1 U1345 ( .B1(n280), .B2(n2089), .C1(n277), .C2(n2057), .A(n958), 
        .ZN(n955) );
  AOI22_X1 U1346 ( .A1(\REGS[23][31] ), .A2(n274), .B1(\REGS[22][31] ), .B2(
        n271), .ZN(n958) );
  OAI221_X1 U1347 ( .B1(n232), .B2(n539), .C1(n229), .C2(n507), .A(n966), .ZN(
        n963) );
  AOI22_X1 U1348 ( .A1(\REGS[7][31] ), .A2(n226), .B1(\REGS[6][31] ), .B2(n223), .ZN(n966) );
  OAI221_X1 U1349 ( .B1(n270), .B2(n2173), .C1(n267), .C2(n2141), .A(n577), 
        .ZN(n562) );
  AOI22_X1 U1350 ( .A1(\REGS[27][11] ), .A2(n264), .B1(\REGS[26][11] ), .B2(
        n261), .ZN(n577) );
  OAI221_X1 U1351 ( .B1(n270), .B2(n2172), .C1(n267), .C2(n2140), .A(n617), 
        .ZN(n612) );
  AOI22_X1 U1352 ( .A1(\REGS[27][12] ), .A2(n264), .B1(\REGS[26][12] ), .B2(
        n261), .ZN(n617) );
  OAI221_X1 U1353 ( .B1(n270), .B2(n2171), .C1(n267), .C2(n2139), .A(n635), 
        .ZN(n630) );
  AOI22_X1 U1354 ( .A1(\REGS[27][13] ), .A2(n264), .B1(\REGS[26][13] ), .B2(
        n261), .ZN(n635) );
  OAI221_X1 U1355 ( .B1(n270), .B2(n2170), .C1(n267), .C2(n2138), .A(n653), 
        .ZN(n648) );
  AOI22_X1 U1356 ( .A1(\REGS[27][14] ), .A2(n264), .B1(\REGS[26][14] ), .B2(
        n261), .ZN(n653) );
  OAI221_X1 U1357 ( .B1(n270), .B2(n2169), .C1(n267), .C2(n2137), .A(n671), 
        .ZN(n666) );
  AOI22_X1 U1358 ( .A1(\REGS[27][15] ), .A2(n264), .B1(\REGS[26][15] ), .B2(
        n261), .ZN(n671) );
  OAI221_X1 U1359 ( .B1(n270), .B2(n2168), .C1(n267), .C2(n2136), .A(n689), 
        .ZN(n684) );
  AOI22_X1 U1360 ( .A1(\REGS[27][16] ), .A2(n264), .B1(\REGS[26][16] ), .B2(
        n261), .ZN(n689) );
  OAI221_X1 U1361 ( .B1(n270), .B2(n2167), .C1(n267), .C2(n2135), .A(n707), 
        .ZN(n702) );
  AOI22_X1 U1362 ( .A1(\REGS[27][17] ), .A2(n264), .B1(\REGS[26][17] ), .B2(
        n261), .ZN(n707) );
  OAI221_X1 U1363 ( .B1(n270), .B2(n2166), .C1(n267), .C2(n2134), .A(n725), 
        .ZN(n720) );
  AOI22_X1 U1364 ( .A1(\REGS[27][18] ), .A2(n264), .B1(\REGS[26][18] ), .B2(
        n261), .ZN(n725) );
  OAI221_X1 U1365 ( .B1(n222), .B2(n1917), .C1(n219), .C2(n1885), .A(n601), 
        .ZN(n586) );
  AOI22_X1 U1366 ( .A1(\REGS[11][11] ), .A2(n216), .B1(\REGS[10][11] ), .B2(
        n213), .ZN(n601) );
  OAI221_X1 U1367 ( .B1(n222), .B2(n1916), .C1(n219), .C2(n1884), .A(n625), 
        .ZN(n620) );
  AOI22_X1 U1368 ( .A1(\REGS[11][12] ), .A2(n216), .B1(\REGS[10][12] ), .B2(
        n213), .ZN(n625) );
  OAI221_X1 U1369 ( .B1(n222), .B2(n1915), .C1(n219), .C2(n1883), .A(n643), 
        .ZN(n638) );
  AOI22_X1 U1370 ( .A1(\REGS[11][13] ), .A2(n216), .B1(\REGS[10][13] ), .B2(
        n213), .ZN(n643) );
  OAI221_X1 U1371 ( .B1(n222), .B2(n1914), .C1(n219), .C2(n1882), .A(n661), 
        .ZN(n656) );
  AOI22_X1 U1372 ( .A1(\REGS[11][14] ), .A2(n216), .B1(\REGS[10][14] ), .B2(
        n213), .ZN(n661) );
  OAI221_X1 U1373 ( .B1(n222), .B2(n1913), .C1(n219), .C2(n1881), .A(n679), 
        .ZN(n674) );
  AOI22_X1 U1374 ( .A1(\REGS[11][15] ), .A2(n216), .B1(\REGS[10][15] ), .B2(
        n213), .ZN(n679) );
  OAI221_X1 U1375 ( .B1(n222), .B2(n1912), .C1(n219), .C2(n1880), .A(n697), 
        .ZN(n692) );
  AOI22_X1 U1376 ( .A1(\REGS[11][16] ), .A2(n216), .B1(\REGS[10][16] ), .B2(
        n213), .ZN(n697) );
  OAI221_X1 U1377 ( .B1(n222), .B2(n1911), .C1(n219), .C2(n1879), .A(n715), 
        .ZN(n710) );
  AOI22_X1 U1378 ( .A1(\REGS[11][17] ), .A2(n216), .B1(\REGS[10][17] ), .B2(
        n213), .ZN(n715) );
  OAI221_X1 U1379 ( .B1(n222), .B2(n1910), .C1(n219), .C2(n1878), .A(n733), 
        .ZN(n728) );
  AOI22_X1 U1380 ( .A1(\REGS[11][18] ), .A2(n216), .B1(\REGS[10][18] ), .B2(
        n213), .ZN(n733) );
  OAI221_X1 U1381 ( .B1(n258), .B2(n2237), .C1(n255), .C2(n2205), .A(n582), 
        .ZN(n561) );
  AOI22_X1 U1382 ( .A1(\REGS[29][11] ), .A2(n252), .B1(\REGS[28][11] ), .B2(
        n249), .ZN(n582) );
  OAI221_X1 U1383 ( .B1(n258), .B2(n2236), .C1(n255), .C2(n2204), .A(n618), 
        .ZN(n611) );
  AOI22_X1 U1384 ( .A1(\REGS[29][12] ), .A2(n252), .B1(\REGS[28][12] ), .B2(
        n249), .ZN(n618) );
  OAI221_X1 U1385 ( .B1(n258), .B2(n2235), .C1(n255), .C2(n2203), .A(n636), 
        .ZN(n629) );
  AOI22_X1 U1386 ( .A1(\REGS[29][13] ), .A2(n252), .B1(\REGS[28][13] ), .B2(
        n249), .ZN(n636) );
  OAI221_X1 U1387 ( .B1(n258), .B2(n2234), .C1(n255), .C2(n2202), .A(n654), 
        .ZN(n647) );
  AOI22_X1 U1388 ( .A1(\REGS[29][14] ), .A2(n252), .B1(\REGS[28][14] ), .B2(
        n249), .ZN(n654) );
  OAI221_X1 U1389 ( .B1(n258), .B2(n2233), .C1(n255), .C2(n2201), .A(n672), 
        .ZN(n665) );
  AOI22_X1 U1390 ( .A1(\REGS[29][15] ), .A2(n252), .B1(\REGS[28][15] ), .B2(
        n249), .ZN(n672) );
  OAI221_X1 U1391 ( .B1(n258), .B2(n2232), .C1(n255), .C2(n2200), .A(n690), 
        .ZN(n683) );
  AOI22_X1 U1392 ( .A1(\REGS[29][16] ), .A2(n252), .B1(\REGS[28][16] ), .B2(
        n249), .ZN(n690) );
  OAI221_X1 U1393 ( .B1(n258), .B2(n2231), .C1(n255), .C2(n2199), .A(n708), 
        .ZN(n701) );
  AOI22_X1 U1394 ( .A1(\REGS[29][17] ), .A2(n252), .B1(\REGS[28][17] ), .B2(
        n249), .ZN(n708) );
  OAI221_X1 U1395 ( .B1(n258), .B2(n2230), .C1(n255), .C2(n2198), .A(n726), 
        .ZN(n719) );
  AOI22_X1 U1396 ( .A1(\REGS[29][18] ), .A2(n252), .B1(\REGS[28][18] ), .B2(
        n249), .ZN(n726) );
  OAI221_X1 U1397 ( .B1(n2159), .B2(n168), .C1(n2127), .C2(n163), .A(n1505), 
        .ZN(n1500) );
  AOI22_X1 U1398 ( .A1(n162), .A2(\REGS[27][25] ), .B1(n159), .B2(
        \REGS[26][25] ), .ZN(n1505) );
  OAI221_X1 U1399 ( .B1(n1903), .B2(n120), .C1(n1871), .C2(n115), .A(n1513), 
        .ZN(n1508) );
  AOI22_X1 U1400 ( .A1(n114), .A2(\REGS[11][25] ), .B1(n111), .B2(
        \REGS[10][25] ), .ZN(n1513) );
  OAI221_X1 U1401 ( .B1(n2158), .B2(n168), .C1(n2126), .C2(n163), .A(n1523), 
        .ZN(n1518) );
  AOI22_X1 U1402 ( .A1(n162), .A2(\REGS[27][26] ), .B1(n159), .B2(
        \REGS[26][26] ), .ZN(n1523) );
  OAI221_X1 U1403 ( .B1(n1902), .B2(n120), .C1(n1870), .C2(n115), .A(n1531), 
        .ZN(n1526) );
  AOI22_X1 U1404 ( .A1(n114), .A2(\REGS[11][26] ), .B1(n111), .B2(
        \REGS[10][26] ), .ZN(n1531) );
  OAI221_X1 U1405 ( .B1(n2157), .B2(n168), .C1(n2125), .C2(n163), .A(n1541), 
        .ZN(n1536) );
  AOI22_X1 U1406 ( .A1(n162), .A2(\REGS[27][27] ), .B1(n159), .B2(
        \REGS[26][27] ), .ZN(n1541) );
  OAI221_X1 U1407 ( .B1(n1901), .B2(n120), .C1(n1869), .C2(n115), .A(n1549), 
        .ZN(n1544) );
  AOI22_X1 U1408 ( .A1(n114), .A2(\REGS[11][27] ), .B1(n111), .B2(
        \REGS[10][27] ), .ZN(n1549) );
  OAI221_X1 U1409 ( .B1(n2156), .B2(n168), .C1(n2124), .C2(n163), .A(n1559), 
        .ZN(n1554) );
  AOI22_X1 U1410 ( .A1(n162), .A2(\REGS[27][28] ), .B1(n159), .B2(
        \REGS[26][28] ), .ZN(n1559) );
  OAI221_X1 U1411 ( .B1(n1900), .B2(n120), .C1(n1868), .C2(n115), .A(n1567), 
        .ZN(n1562) );
  AOI22_X1 U1412 ( .A1(n114), .A2(\REGS[11][28] ), .B1(n111), .B2(
        \REGS[10][28] ), .ZN(n1567) );
  OAI221_X1 U1413 ( .B1(n2155), .B2(n168), .C1(n2123), .C2(n163), .A(n1577), 
        .ZN(n1572) );
  AOI22_X1 U1414 ( .A1(n162), .A2(\REGS[27][29] ), .B1(n159), .B2(
        \REGS[26][29] ), .ZN(n1577) );
  OAI221_X1 U1415 ( .B1(n1899), .B2(n120), .C1(n1867), .C2(n115), .A(n1585), 
        .ZN(n1580) );
  AOI22_X1 U1416 ( .A1(n114), .A2(\REGS[11][29] ), .B1(n111), .B2(
        \REGS[10][29] ), .ZN(n1585) );
  OAI221_X1 U1417 ( .B1(n2154), .B2(n168), .C1(n2122), .C2(n163), .A(n1595), 
        .ZN(n1590) );
  AOI22_X1 U1418 ( .A1(n162), .A2(\REGS[27][30] ), .B1(n159), .B2(
        \REGS[26][30] ), .ZN(n1595) );
  OAI221_X1 U1419 ( .B1(n1898), .B2(n120), .C1(n1866), .C2(n115), .A(n1603), 
        .ZN(n1598) );
  AOI22_X1 U1420 ( .A1(n114), .A2(\REGS[11][30] ), .B1(n111), .B2(
        \REGS[10][30] ), .ZN(n1603) );
  OAI221_X1 U1421 ( .B1(n2153), .B2(n168), .C1(n2121), .C2(n163), .A(n1620), 
        .ZN(n1608) );
  AOI22_X1 U1422 ( .A1(n162), .A2(\REGS[27][31] ), .B1(n159), .B2(
        \REGS[26][31] ), .ZN(n1620) );
  OAI221_X1 U1423 ( .B1(n1897), .B2(n120), .C1(n1865), .C2(n115), .A(n1634), 
        .ZN(n1626) );
  AOI22_X1 U1424 ( .A1(n114), .A2(\REGS[11][31] ), .B1(n111), .B2(
        \REGS[10][31] ), .ZN(n1634) );
  OAI221_X1 U1425 ( .B1(n2223), .B2(n156), .C1(n2191), .C2(n151), .A(n1506), 
        .ZN(n1499) );
  AOI22_X1 U1426 ( .A1(n150), .A2(\REGS[29][25] ), .B1(n147), .B2(
        \REGS[28][25] ), .ZN(n1506) );
  OAI221_X1 U1427 ( .B1(n2222), .B2(n156), .C1(n2190), .C2(n151), .A(n1524), 
        .ZN(n1517) );
  AOI22_X1 U1428 ( .A1(n150), .A2(\REGS[29][26] ), .B1(n147), .B2(
        \REGS[28][26] ), .ZN(n1524) );
  OAI221_X1 U1429 ( .B1(n2221), .B2(n156), .C1(n2189), .C2(n151), .A(n1542), 
        .ZN(n1535) );
  AOI22_X1 U1430 ( .A1(n150), .A2(\REGS[29][27] ), .B1(n147), .B2(
        \REGS[28][27] ), .ZN(n1542) );
  OAI221_X1 U1431 ( .B1(n2220), .B2(n156), .C1(n2188), .C2(n151), .A(n1560), 
        .ZN(n1553) );
  AOI22_X1 U1432 ( .A1(n150), .A2(\REGS[29][28] ), .B1(n147), .B2(
        \REGS[28][28] ), .ZN(n1560) );
  OAI221_X1 U1433 ( .B1(n2219), .B2(n156), .C1(n2187), .C2(n151), .A(n1578), 
        .ZN(n1571) );
  AOI22_X1 U1434 ( .A1(n150), .A2(\REGS[29][29] ), .B1(n147), .B2(
        \REGS[28][29] ), .ZN(n1578) );
  OAI221_X1 U1435 ( .B1(n2218), .B2(n156), .C1(n2186), .C2(n151), .A(n1596), 
        .ZN(n1589) );
  AOI22_X1 U1436 ( .A1(n150), .A2(\REGS[29][30] ), .B1(n147), .B2(
        \REGS[28][30] ), .ZN(n1596) );
  OAI221_X1 U1437 ( .B1(n2217), .B2(n156), .C1(n2185), .C2(n151), .A(n1623), 
        .ZN(n1607) );
  AOI22_X1 U1438 ( .A1(n150), .A2(\REGS[29][31] ), .B1(n147), .B2(
        \REGS[28][31] ), .ZN(n1623) );
  OAI221_X1 U1439 ( .B1(n268), .B2(n2184), .C1(n265), .C2(n2152), .A(n1647), 
        .ZN(n1642) );
  AOI22_X1 U1440 ( .A1(\REGS[27][0] ), .A2(n262), .B1(\REGS[26][0] ), .B2(n259), .ZN(n1647) );
  OAI221_X1 U1441 ( .B1(n220), .B2(n1928), .C1(n217), .C2(n1896), .A(n1655), 
        .ZN(n1650) );
  AOI22_X1 U1442 ( .A1(\REGS[11][0] ), .A2(n214), .B1(\REGS[10][0] ), .B2(n211), .ZN(n1655) );
  OAI221_X1 U1443 ( .B1(n166), .B2(n2184), .C1(n165), .C2(n2152), .A(n1033), 
        .ZN(n1018) );
  AOI22_X1 U1444 ( .A1(\REGS[27][0] ), .A2(n160), .B1(\REGS[26][0] ), .B2(n157), .ZN(n1033) );
  OAI221_X1 U1445 ( .B1(n118), .B2(n1928), .C1(n117), .C2(n1896), .A(n1057), 
        .ZN(n1042) );
  AOI22_X1 U1446 ( .A1(\REGS[11][0] ), .A2(n112), .B1(\REGS[10][0] ), .B2(n109), .ZN(n1057) );
  OAI221_X1 U1447 ( .B1(n268), .B2(n2183), .C1(n265), .C2(n2151), .A(n1665), 
        .ZN(n1660) );
  AOI22_X1 U1448 ( .A1(\REGS[27][1] ), .A2(n262), .B1(\REGS[26][1] ), .B2(n259), .ZN(n1665) );
  OAI221_X1 U1449 ( .B1(n220), .B2(n1927), .C1(n217), .C2(n1895), .A(n1673), 
        .ZN(n1668) );
  AOI22_X1 U1450 ( .A1(\REGS[11][1] ), .A2(n214), .B1(\REGS[10][1] ), .B2(n211), .ZN(n1673) );
  OAI221_X1 U1451 ( .B1(n166), .B2(n2183), .C1(n165), .C2(n2151), .A(n1073), 
        .ZN(n1068) );
  AOI22_X1 U1452 ( .A1(\REGS[27][1] ), .A2(n160), .B1(\REGS[26][1] ), .B2(n157), .ZN(n1073) );
  OAI221_X1 U1453 ( .B1(n118), .B2(n1927), .C1(n117), .C2(n1895), .A(n1081), 
        .ZN(n1076) );
  AOI22_X1 U1454 ( .A1(\REGS[11][1] ), .A2(n112), .B1(\REGS[10][1] ), .B2(n109), .ZN(n1081) );
  OAI221_X1 U1455 ( .B1(n268), .B2(n2182), .C1(n265), .C2(n2150), .A(n1683), 
        .ZN(n1678) );
  AOI22_X1 U1456 ( .A1(\REGS[27][2] ), .A2(n262), .B1(\REGS[26][2] ), .B2(n259), .ZN(n1683) );
  OAI221_X1 U1457 ( .B1(n220), .B2(n1926), .C1(n217), .C2(n1894), .A(n1691), 
        .ZN(n1686) );
  AOI22_X1 U1458 ( .A1(\REGS[11][2] ), .A2(n214), .B1(\REGS[10][2] ), .B2(n211), .ZN(n1691) );
  OAI221_X1 U1459 ( .B1(n166), .B2(n2182), .C1(n165), .C2(n2150), .A(n1091), 
        .ZN(n1086) );
  AOI22_X1 U1460 ( .A1(\REGS[27][2] ), .A2(n160), .B1(\REGS[26][2] ), .B2(n157), .ZN(n1091) );
  OAI221_X1 U1461 ( .B1(n118), .B2(n1926), .C1(n117), .C2(n1894), .A(n1099), 
        .ZN(n1094) );
  AOI22_X1 U1462 ( .A1(\REGS[11][2] ), .A2(n112), .B1(\REGS[10][2] ), .B2(n109), .ZN(n1099) );
  OAI221_X1 U1463 ( .B1(n268), .B2(n2181), .C1(n265), .C2(n2149), .A(n1701), 
        .ZN(n1696) );
  AOI22_X1 U1464 ( .A1(\REGS[27][3] ), .A2(n262), .B1(\REGS[26][3] ), .B2(n259), .ZN(n1701) );
  OAI221_X1 U1465 ( .B1(n220), .B2(n1925), .C1(n217), .C2(n1893), .A(n1709), 
        .ZN(n1704) );
  AOI22_X1 U1466 ( .A1(\REGS[11][3] ), .A2(n214), .B1(\REGS[10][3] ), .B2(n211), .ZN(n1709) );
  OAI221_X1 U1467 ( .B1(n166), .B2(n2181), .C1(n165), .C2(n2149), .A(n1109), 
        .ZN(n1104) );
  AOI22_X1 U1468 ( .A1(\REGS[27][3] ), .A2(n160), .B1(\REGS[26][3] ), .B2(n157), .ZN(n1109) );
  OAI221_X1 U1469 ( .B1(n118), .B2(n1925), .C1(n117), .C2(n1893), .A(n1117), 
        .ZN(n1112) );
  AOI22_X1 U1470 ( .A1(\REGS[11][3] ), .A2(n112), .B1(\REGS[10][3] ), .B2(n109), .ZN(n1117) );
  OAI221_X1 U1471 ( .B1(n268), .B2(n2180), .C1(n265), .C2(n2148), .A(n1719), 
        .ZN(n1714) );
  AOI22_X1 U1472 ( .A1(\REGS[27][4] ), .A2(n262), .B1(\REGS[26][4] ), .B2(n259), .ZN(n1719) );
  OAI221_X1 U1473 ( .B1(n220), .B2(n1924), .C1(n217), .C2(n1892), .A(n1727), 
        .ZN(n1722) );
  AOI22_X1 U1474 ( .A1(\REGS[11][4] ), .A2(n214), .B1(\REGS[10][4] ), .B2(n211), .ZN(n1727) );
  OAI221_X1 U1475 ( .B1(n166), .B2(n2180), .C1(n165), .C2(n2148), .A(n1127), 
        .ZN(n1122) );
  AOI22_X1 U1476 ( .A1(\REGS[27][4] ), .A2(n160), .B1(\REGS[26][4] ), .B2(n157), .ZN(n1127) );
  OAI221_X1 U1477 ( .B1(n118), .B2(n1924), .C1(n117), .C2(n1892), .A(n1135), 
        .ZN(n1130) );
  AOI22_X1 U1478 ( .A1(\REGS[11][4] ), .A2(n112), .B1(\REGS[10][4] ), .B2(n109), .ZN(n1135) );
  OAI221_X1 U1479 ( .B1(n268), .B2(n2179), .C1(n265), .C2(n2147), .A(n1737), 
        .ZN(n1732) );
  AOI22_X1 U1480 ( .A1(\REGS[27][5] ), .A2(n262), .B1(\REGS[26][5] ), .B2(n259), .ZN(n1737) );
  OAI221_X1 U1481 ( .B1(n220), .B2(n1923), .C1(n217), .C2(n1891), .A(n1745), 
        .ZN(n1740) );
  AOI22_X1 U1482 ( .A1(\REGS[11][5] ), .A2(n214), .B1(\REGS[10][5] ), .B2(n211), .ZN(n1745) );
  OAI221_X1 U1483 ( .B1(n166), .B2(n2179), .C1(n165), .C2(n2147), .A(n1145), 
        .ZN(n1140) );
  AOI22_X1 U1484 ( .A1(\REGS[27][5] ), .A2(n160), .B1(\REGS[26][5] ), .B2(n157), .ZN(n1145) );
  OAI221_X1 U1485 ( .B1(n118), .B2(n1923), .C1(n117), .C2(n1891), .A(n1153), 
        .ZN(n1148) );
  AOI22_X1 U1486 ( .A1(\REGS[11][5] ), .A2(n112), .B1(\REGS[10][5] ), .B2(n109), .ZN(n1153) );
  OAI221_X1 U1487 ( .B1(n268), .B2(n2178), .C1(n265), .C2(n2146), .A(n1755), 
        .ZN(n1750) );
  AOI22_X1 U1488 ( .A1(\REGS[27][6] ), .A2(n262), .B1(\REGS[26][6] ), .B2(n259), .ZN(n1755) );
  OAI221_X1 U1489 ( .B1(n220), .B2(n1922), .C1(n217), .C2(n1890), .A(n1763), 
        .ZN(n1758) );
  AOI22_X1 U1490 ( .A1(\REGS[11][6] ), .A2(n214), .B1(\REGS[10][6] ), .B2(n211), .ZN(n1763) );
  OAI221_X1 U1491 ( .B1(n166), .B2(n2178), .C1(n165), .C2(n2146), .A(n1163), 
        .ZN(n1158) );
  AOI22_X1 U1492 ( .A1(\REGS[27][6] ), .A2(n160), .B1(\REGS[26][6] ), .B2(n157), .ZN(n1163) );
  OAI221_X1 U1493 ( .B1(n118), .B2(n1922), .C1(n117), .C2(n1890), .A(n1171), 
        .ZN(n1166) );
  AOI22_X1 U1494 ( .A1(\REGS[11][6] ), .A2(n112), .B1(\REGS[10][6] ), .B2(n109), .ZN(n1171) );
  OAI221_X1 U1495 ( .B1(n268), .B2(n2177), .C1(n265), .C2(n2145), .A(n1773), 
        .ZN(n1768) );
  AOI22_X1 U1496 ( .A1(\REGS[27][7] ), .A2(n262), .B1(\REGS[26][7] ), .B2(n259), .ZN(n1773) );
  OAI221_X1 U1497 ( .B1(n220), .B2(n1921), .C1(n217), .C2(n1889), .A(n1781), 
        .ZN(n1776) );
  AOI22_X1 U1498 ( .A1(\REGS[11][7] ), .A2(n214), .B1(\REGS[10][7] ), .B2(n211), .ZN(n1781) );
  OAI221_X1 U1499 ( .B1(n166), .B2(n2177), .C1(n165), .C2(n2145), .A(n1181), 
        .ZN(n1176) );
  AOI22_X1 U1500 ( .A1(\REGS[27][7] ), .A2(n160), .B1(\REGS[26][7] ), .B2(n157), .ZN(n1181) );
  OAI221_X1 U1501 ( .B1(n118), .B2(n1921), .C1(n117), .C2(n1889), .A(n1189), 
        .ZN(n1184) );
  AOI22_X1 U1502 ( .A1(\REGS[11][7] ), .A2(n112), .B1(\REGS[10][7] ), .B2(n109), .ZN(n1189) );
  OAI221_X1 U1503 ( .B1(n268), .B2(n2176), .C1(n265), .C2(n2144), .A(n1791), 
        .ZN(n1786) );
  AOI22_X1 U1504 ( .A1(\REGS[27][8] ), .A2(n262), .B1(\REGS[26][8] ), .B2(n259), .ZN(n1791) );
  OAI221_X1 U1505 ( .B1(n220), .B2(n1920), .C1(n217), .C2(n1888), .A(n1799), 
        .ZN(n1794) );
  AOI22_X1 U1506 ( .A1(\REGS[11][8] ), .A2(n214), .B1(\REGS[10][8] ), .B2(n211), .ZN(n1799) );
  OAI221_X1 U1507 ( .B1(n166), .B2(n2176), .C1(n164), .C2(n2144), .A(n1199), 
        .ZN(n1194) );
  AOI22_X1 U1508 ( .A1(\REGS[27][8] ), .A2(n160), .B1(\REGS[26][8] ), .B2(n157), .ZN(n1199) );
  OAI221_X1 U1509 ( .B1(n118), .B2(n1920), .C1(n116), .C2(n1888), .A(n1207), 
        .ZN(n1202) );
  AOI22_X1 U1510 ( .A1(\REGS[11][8] ), .A2(n112), .B1(\REGS[10][8] ), .B2(n109), .ZN(n1207) );
  OAI221_X1 U1511 ( .B1(n268), .B2(n2175), .C1(n265), .C2(n2143), .A(n1809), 
        .ZN(n1804) );
  AOI22_X1 U1512 ( .A1(\REGS[27][9] ), .A2(n262), .B1(\REGS[26][9] ), .B2(n259), .ZN(n1809) );
  OAI221_X1 U1513 ( .B1(n220), .B2(n1919), .C1(n217), .C2(n1887), .A(n1817), 
        .ZN(n1812) );
  AOI22_X1 U1514 ( .A1(\REGS[11][9] ), .A2(n214), .B1(\REGS[10][9] ), .B2(n211), .ZN(n1817) );
  OAI221_X1 U1515 ( .B1(n166), .B2(n2175), .C1(n164), .C2(n2143), .A(n1217), 
        .ZN(n1212) );
  AOI22_X1 U1516 ( .A1(\REGS[27][9] ), .A2(n160), .B1(\REGS[26][9] ), .B2(n157), .ZN(n1217) );
  OAI221_X1 U1517 ( .B1(n118), .B2(n1919), .C1(n116), .C2(n1887), .A(n1225), 
        .ZN(n1220) );
  AOI22_X1 U1518 ( .A1(\REGS[11][9] ), .A2(n112), .B1(\REGS[10][9] ), .B2(n109), .ZN(n1225) );
  OAI221_X1 U1519 ( .B1(n268), .B2(n2174), .C1(n265), .C2(n2142), .A(n1834), 
        .ZN(n1822) );
  AOI22_X1 U1520 ( .A1(\REGS[27][10] ), .A2(n262), .B1(\REGS[26][10] ), .B2(
        n259), .ZN(n1834) );
  OAI221_X1 U1521 ( .B1(n220), .B2(n1918), .C1(n217), .C2(n1886), .A(n1848), 
        .ZN(n1840) );
  AOI22_X1 U1522 ( .A1(\REGS[11][10] ), .A2(n214), .B1(\REGS[10][10] ), .B2(
        n211), .ZN(n1848) );
  OAI221_X1 U1523 ( .B1(n166), .B2(n2174), .C1(n164), .C2(n2142), .A(n1235), 
        .ZN(n1230) );
  AOI22_X1 U1524 ( .A1(\REGS[27][10] ), .A2(n160), .B1(\REGS[26][10] ), .B2(
        n157), .ZN(n1235) );
  OAI221_X1 U1525 ( .B1(n118), .B2(n1918), .C1(n116), .C2(n1886), .A(n1243), 
        .ZN(n1238) );
  AOI22_X1 U1526 ( .A1(\REGS[11][10] ), .A2(n112), .B1(\REGS[10][10] ), .B2(
        n109), .ZN(n1243) );
  OAI221_X1 U1527 ( .B1(n2173), .B2(n166), .C1(n2141), .C2(n164), .A(n1253), 
        .ZN(n1248) );
  AOI22_X1 U1528 ( .A1(n160), .A2(\REGS[27][11] ), .B1(n157), .B2(
        \REGS[26][11] ), .ZN(n1253) );
  OAI221_X1 U1529 ( .B1(n1917), .B2(n118), .C1(n1885), .C2(n116), .A(n1261), 
        .ZN(n1256) );
  AOI22_X1 U1530 ( .A1(n112), .A2(\REGS[11][11] ), .B1(n109), .B2(
        \REGS[10][11] ), .ZN(n1261) );
  OAI221_X1 U1531 ( .B1(n2172), .B2(n167), .C1(n2140), .C2(n164), .A(n1271), 
        .ZN(n1266) );
  AOI22_X1 U1532 ( .A1(n161), .A2(\REGS[27][12] ), .B1(n158), .B2(
        \REGS[26][12] ), .ZN(n1271) );
  OAI221_X1 U1533 ( .B1(n1916), .B2(n119), .C1(n1884), .C2(n116), .A(n1279), 
        .ZN(n1274) );
  AOI22_X1 U1534 ( .A1(n113), .A2(\REGS[11][12] ), .B1(n110), .B2(
        \REGS[10][12] ), .ZN(n1279) );
  OAI221_X1 U1535 ( .B1(n2171), .B2(n167), .C1(n2139), .C2(n164), .A(n1289), 
        .ZN(n1284) );
  AOI22_X1 U1536 ( .A1(n161), .A2(\REGS[27][13] ), .B1(n158), .B2(
        \REGS[26][13] ), .ZN(n1289) );
  OAI221_X1 U1537 ( .B1(n1915), .B2(n119), .C1(n1883), .C2(n116), .A(n1297), 
        .ZN(n1292) );
  AOI22_X1 U1538 ( .A1(n113), .A2(\REGS[11][13] ), .B1(n110), .B2(
        \REGS[10][13] ), .ZN(n1297) );
  OAI221_X1 U1539 ( .B1(n2170), .B2(n167), .C1(n2138), .C2(n164), .A(n1307), 
        .ZN(n1302) );
  AOI22_X1 U1540 ( .A1(n161), .A2(\REGS[27][14] ), .B1(n158), .B2(
        \REGS[26][14] ), .ZN(n1307) );
  OAI221_X1 U1541 ( .B1(n1914), .B2(n119), .C1(n1882), .C2(n116), .A(n1315), 
        .ZN(n1310) );
  AOI22_X1 U1542 ( .A1(n113), .A2(\REGS[11][14] ), .B1(n110), .B2(
        \REGS[10][14] ), .ZN(n1315) );
  OAI221_X1 U1543 ( .B1(n2169), .B2(n167), .C1(n2137), .C2(n164), .A(n1325), 
        .ZN(n1320) );
  AOI22_X1 U1544 ( .A1(n161), .A2(\REGS[27][15] ), .B1(n158), .B2(
        \REGS[26][15] ), .ZN(n1325) );
  OAI221_X1 U1545 ( .B1(n1913), .B2(n119), .C1(n1881), .C2(n116), .A(n1333), 
        .ZN(n1328) );
  AOI22_X1 U1546 ( .A1(n113), .A2(\REGS[11][15] ), .B1(n110), .B2(
        \REGS[10][15] ), .ZN(n1333) );
  OAI221_X1 U1547 ( .B1(n2168), .B2(n167), .C1(n2136), .C2(n164), .A(n1343), 
        .ZN(n1338) );
  AOI22_X1 U1548 ( .A1(n161), .A2(\REGS[27][16] ), .B1(n158), .B2(
        \REGS[26][16] ), .ZN(n1343) );
  OAI221_X1 U1549 ( .B1(n1912), .B2(n119), .C1(n1880), .C2(n116), .A(n1351), 
        .ZN(n1346) );
  AOI22_X1 U1550 ( .A1(n113), .A2(\REGS[11][16] ), .B1(n110), .B2(
        \REGS[10][16] ), .ZN(n1351) );
  OAI221_X1 U1551 ( .B1(n2167), .B2(n167), .C1(n2135), .C2(n164), .A(n1361), 
        .ZN(n1356) );
  AOI22_X1 U1552 ( .A1(n161), .A2(\REGS[27][17] ), .B1(n158), .B2(
        \REGS[26][17] ), .ZN(n1361) );
  OAI221_X1 U1553 ( .B1(n1911), .B2(n119), .C1(n1879), .C2(n116), .A(n1369), 
        .ZN(n1364) );
  AOI22_X1 U1554 ( .A1(n113), .A2(\REGS[11][17] ), .B1(n110), .B2(
        \REGS[10][17] ), .ZN(n1369) );
  OAI221_X1 U1555 ( .B1(n2166), .B2(n167), .C1(n2134), .C2(n164), .A(n1379), 
        .ZN(n1374) );
  AOI22_X1 U1556 ( .A1(n161), .A2(\REGS[27][18] ), .B1(n158), .B2(
        \REGS[26][18] ), .ZN(n1379) );
  OAI221_X1 U1557 ( .B1(n1910), .B2(n119), .C1(n1878), .C2(n116), .A(n1387), 
        .ZN(n1382) );
  AOI22_X1 U1558 ( .A1(n113), .A2(\REGS[11][18] ), .B1(n110), .B2(
        \REGS[10][18] ), .ZN(n1387) );
  OAI221_X1 U1559 ( .B1(n2165), .B2(n167), .C1(n2133), .C2(n164), .A(n1397), 
        .ZN(n1392) );
  AOI22_X1 U1560 ( .A1(n161), .A2(\REGS[27][19] ), .B1(n158), .B2(
        \REGS[26][19] ), .ZN(n1397) );
  OAI221_X1 U1561 ( .B1(n1909), .B2(n119), .C1(n1877), .C2(n116), .A(n1405), 
        .ZN(n1400) );
  AOI22_X1 U1562 ( .A1(n113), .A2(\REGS[11][19] ), .B1(n110), .B2(
        \REGS[10][19] ), .ZN(n1405) );
  OAI221_X1 U1563 ( .B1(n269), .B2(n2165), .C1(n266), .C2(n2133), .A(n743), 
        .ZN(n738) );
  AOI22_X1 U1564 ( .A1(\REGS[27][19] ), .A2(n263), .B1(\REGS[26][19] ), .B2(
        n260), .ZN(n743) );
  OAI221_X1 U1565 ( .B1(n221), .B2(n1909), .C1(n218), .C2(n1877), .A(n751), 
        .ZN(n746) );
  AOI22_X1 U1566 ( .A1(\REGS[11][19] ), .A2(n215), .B1(\REGS[10][19] ), .B2(
        n212), .ZN(n751) );
  OAI221_X1 U1567 ( .B1(n2164), .B2(n167), .C1(n2132), .C2(n163), .A(n1415), 
        .ZN(n1410) );
  AOI22_X1 U1568 ( .A1(n161), .A2(\REGS[27][20] ), .B1(n158), .B2(
        \REGS[26][20] ), .ZN(n1415) );
  OAI221_X1 U1569 ( .B1(n1908), .B2(n119), .C1(n1876), .C2(n115), .A(n1423), 
        .ZN(n1418) );
  AOI22_X1 U1570 ( .A1(n113), .A2(\REGS[11][20] ), .B1(n110), .B2(
        \REGS[10][20] ), .ZN(n1423) );
  OAI221_X1 U1571 ( .B1(n269), .B2(n2164), .C1(n266), .C2(n2132), .A(n761), 
        .ZN(n756) );
  AOI22_X1 U1572 ( .A1(\REGS[27][20] ), .A2(n263), .B1(\REGS[26][20] ), .B2(
        n260), .ZN(n761) );
  OAI221_X1 U1573 ( .B1(n221), .B2(n1908), .C1(n218), .C2(n1876), .A(n769), 
        .ZN(n764) );
  AOI22_X1 U1574 ( .A1(\REGS[11][20] ), .A2(n215), .B1(\REGS[10][20] ), .B2(
        n212), .ZN(n769) );
  OAI221_X1 U1575 ( .B1(n2163), .B2(n167), .C1(n2131), .C2(n163), .A(n1433), 
        .ZN(n1428) );
  AOI22_X1 U1576 ( .A1(n161), .A2(\REGS[27][21] ), .B1(n158), .B2(
        \REGS[26][21] ), .ZN(n1433) );
  OAI221_X1 U1577 ( .B1(n1907), .B2(n119), .C1(n1875), .C2(n115), .A(n1441), 
        .ZN(n1436) );
  AOI22_X1 U1578 ( .A1(n113), .A2(\REGS[11][21] ), .B1(n110), .B2(
        \REGS[10][21] ), .ZN(n1441) );
  OAI221_X1 U1579 ( .B1(n269), .B2(n2163), .C1(n266), .C2(n2131), .A(n779), 
        .ZN(n774) );
  AOI22_X1 U1580 ( .A1(\REGS[27][21] ), .A2(n263), .B1(\REGS[26][21] ), .B2(
        n260), .ZN(n779) );
  OAI221_X1 U1581 ( .B1(n221), .B2(n1907), .C1(n218), .C2(n1875), .A(n787), 
        .ZN(n782) );
  AOI22_X1 U1582 ( .A1(\REGS[11][21] ), .A2(n215), .B1(\REGS[10][21] ), .B2(
        n212), .ZN(n787) );
  OAI221_X1 U1583 ( .B1(n2162), .B2(n167), .C1(n2130), .C2(n163), .A(n1451), 
        .ZN(n1446) );
  AOI22_X1 U1584 ( .A1(n161), .A2(\REGS[27][22] ), .B1(n158), .B2(
        \REGS[26][22] ), .ZN(n1451) );
  OAI221_X1 U1585 ( .B1(n1906), .B2(n119), .C1(n1874), .C2(n115), .A(n1459), 
        .ZN(n1454) );
  AOI22_X1 U1586 ( .A1(n113), .A2(\REGS[11][22] ), .B1(n110), .B2(
        \REGS[10][22] ), .ZN(n1459) );
  OAI221_X1 U1587 ( .B1(n269), .B2(n2162), .C1(n266), .C2(n2130), .A(n797), 
        .ZN(n792) );
  AOI22_X1 U1588 ( .A1(\REGS[27][22] ), .A2(n263), .B1(\REGS[26][22] ), .B2(
        n260), .ZN(n797) );
  OAI221_X1 U1589 ( .B1(n221), .B2(n1906), .C1(n218), .C2(n1874), .A(n805), 
        .ZN(n800) );
  AOI22_X1 U1590 ( .A1(\REGS[11][22] ), .A2(n215), .B1(\REGS[10][22] ), .B2(
        n212), .ZN(n805) );
  OAI221_X1 U1591 ( .B1(n2161), .B2(n167), .C1(n2129), .C2(n163), .A(n1469), 
        .ZN(n1464) );
  AOI22_X1 U1592 ( .A1(n161), .A2(\REGS[27][23] ), .B1(n158), .B2(
        \REGS[26][23] ), .ZN(n1469) );
  OAI221_X1 U1593 ( .B1(n1905), .B2(n119), .C1(n1873), .C2(n115), .A(n1477), 
        .ZN(n1472) );
  AOI22_X1 U1594 ( .A1(n113), .A2(\REGS[11][23] ), .B1(n110), .B2(
        \REGS[10][23] ), .ZN(n1477) );
  OAI221_X1 U1595 ( .B1(n269), .B2(n2161), .C1(n266), .C2(n2129), .A(n815), 
        .ZN(n810) );
  AOI22_X1 U1596 ( .A1(\REGS[27][23] ), .A2(n263), .B1(\REGS[26][23] ), .B2(
        n260), .ZN(n815) );
  OAI221_X1 U1597 ( .B1(n221), .B2(n1905), .C1(n218), .C2(n1873), .A(n823), 
        .ZN(n818) );
  AOI22_X1 U1598 ( .A1(\REGS[11][23] ), .A2(n215), .B1(\REGS[10][23] ), .B2(
        n212), .ZN(n823) );
  OAI221_X1 U1599 ( .B1(n2160), .B2(n167), .C1(n2128), .C2(n163), .A(n1487), 
        .ZN(n1482) );
  AOI22_X1 U1600 ( .A1(n161), .A2(\REGS[27][24] ), .B1(n158), .B2(
        \REGS[26][24] ), .ZN(n1487) );
  OAI221_X1 U1601 ( .B1(n1904), .B2(n119), .C1(n1872), .C2(n115), .A(n1495), 
        .ZN(n1490) );
  AOI22_X1 U1602 ( .A1(n113), .A2(\REGS[11][24] ), .B1(n110), .B2(
        \REGS[10][24] ), .ZN(n1495) );
  OAI221_X1 U1603 ( .B1(n269), .B2(n2160), .C1(n266), .C2(n2128), .A(n833), 
        .ZN(n828) );
  AOI22_X1 U1604 ( .A1(\REGS[27][24] ), .A2(n263), .B1(\REGS[26][24] ), .B2(
        n260), .ZN(n833) );
  OAI221_X1 U1605 ( .B1(n221), .B2(n1904), .C1(n218), .C2(n1872), .A(n841), 
        .ZN(n836) );
  AOI22_X1 U1606 ( .A1(\REGS[11][24] ), .A2(n215), .B1(\REGS[10][24] ), .B2(
        n212), .ZN(n841) );
  OAI221_X1 U1607 ( .B1(n269), .B2(n2159), .C1(n266), .C2(n2127), .A(n851), 
        .ZN(n846) );
  AOI22_X1 U1608 ( .A1(\REGS[27][25] ), .A2(n263), .B1(\REGS[26][25] ), .B2(
        n260), .ZN(n851) );
  OAI221_X1 U1609 ( .B1(n221), .B2(n1903), .C1(n218), .C2(n1871), .A(n859), 
        .ZN(n854) );
  AOI22_X1 U1610 ( .A1(\REGS[11][25] ), .A2(n215), .B1(\REGS[10][25] ), .B2(
        n212), .ZN(n859) );
  OAI221_X1 U1611 ( .B1(n269), .B2(n2158), .C1(n266), .C2(n2126), .A(n869), 
        .ZN(n864) );
  AOI22_X1 U1612 ( .A1(\REGS[27][26] ), .A2(n263), .B1(\REGS[26][26] ), .B2(
        n260), .ZN(n869) );
  OAI221_X1 U1613 ( .B1(n221), .B2(n1902), .C1(n218), .C2(n1870), .A(n877), 
        .ZN(n872) );
  AOI22_X1 U1614 ( .A1(\REGS[11][26] ), .A2(n215), .B1(\REGS[10][26] ), .B2(
        n212), .ZN(n877) );
  OAI221_X1 U1615 ( .B1(n269), .B2(n2157), .C1(n266), .C2(n2125), .A(n887), 
        .ZN(n882) );
  AOI22_X1 U1616 ( .A1(\REGS[27][27] ), .A2(n263), .B1(\REGS[26][27] ), .B2(
        n260), .ZN(n887) );
  OAI221_X1 U1617 ( .B1(n221), .B2(n1901), .C1(n218), .C2(n1869), .A(n895), 
        .ZN(n890) );
  AOI22_X1 U1618 ( .A1(\REGS[11][27] ), .A2(n215), .B1(\REGS[10][27] ), .B2(
        n212), .ZN(n895) );
  OAI221_X1 U1619 ( .B1(n269), .B2(n2156), .C1(n266), .C2(n2124), .A(n905), 
        .ZN(n900) );
  AOI22_X1 U1620 ( .A1(\REGS[27][28] ), .A2(n263), .B1(\REGS[26][28] ), .B2(
        n260), .ZN(n905) );
  OAI221_X1 U1621 ( .B1(n221), .B2(n1900), .C1(n218), .C2(n1868), .A(n913), 
        .ZN(n908) );
  AOI22_X1 U1622 ( .A1(\REGS[11][28] ), .A2(n215), .B1(\REGS[10][28] ), .B2(
        n212), .ZN(n913) );
  OAI221_X1 U1623 ( .B1(n269), .B2(n2155), .C1(n266), .C2(n2123), .A(n923), 
        .ZN(n918) );
  AOI22_X1 U1624 ( .A1(\REGS[27][29] ), .A2(n263), .B1(\REGS[26][29] ), .B2(
        n260), .ZN(n923) );
  OAI221_X1 U1625 ( .B1(n221), .B2(n1899), .C1(n218), .C2(n1867), .A(n931), 
        .ZN(n926) );
  AOI22_X1 U1626 ( .A1(\REGS[11][29] ), .A2(n215), .B1(\REGS[10][29] ), .B2(
        n212), .ZN(n931) );
  OAI221_X1 U1627 ( .B1(n269), .B2(n2154), .C1(n266), .C2(n2122), .A(n941), 
        .ZN(n936) );
  AOI22_X1 U1628 ( .A1(\REGS[27][30] ), .A2(n263), .B1(\REGS[26][30] ), .B2(
        n260), .ZN(n941) );
  OAI221_X1 U1629 ( .B1(n221), .B2(n1898), .C1(n218), .C2(n1866), .A(n949), 
        .ZN(n944) );
  AOI22_X1 U1630 ( .A1(\REGS[11][30] ), .A2(n215), .B1(\REGS[10][30] ), .B2(
        n212), .ZN(n949) );
  OAI221_X1 U1631 ( .B1(n268), .B2(n2153), .C1(n265), .C2(n2121), .A(n959), 
        .ZN(n954) );
  AOI22_X1 U1632 ( .A1(\REGS[27][31] ), .A2(n262), .B1(\REGS[26][31] ), .B2(
        n259), .ZN(n959) );
  OAI221_X1 U1633 ( .B1(n220), .B2(n1897), .C1(n217), .C2(n1865), .A(n967), 
        .ZN(n962) );
  AOI22_X1 U1634 ( .A1(\REGS[11][31] ), .A2(n214), .B1(\REGS[10][31] ), .B2(
        n211), .ZN(n967) );
  OAI221_X1 U1635 ( .B1(n256), .B2(n2248), .C1(n253), .C2(n2216), .A(n1648), 
        .ZN(n1641) );
  AOI22_X1 U1636 ( .A1(\REGS[29][0] ), .A2(n250), .B1(\REGS[28][0] ), .B2(n247), .ZN(n1648) );
  OAI221_X1 U1637 ( .B1(n154), .B2(n2248), .C1(n153), .C2(n2216), .A(n1038), 
        .ZN(n1017) );
  AOI22_X1 U1638 ( .A1(\REGS[29][0] ), .A2(n148), .B1(\REGS[28][0] ), .B2(n145), .ZN(n1038) );
  OAI221_X1 U1639 ( .B1(n256), .B2(n2247), .C1(n253), .C2(n2215), .A(n1666), 
        .ZN(n1659) );
  AOI22_X1 U1640 ( .A1(\REGS[29][1] ), .A2(n250), .B1(\REGS[28][1] ), .B2(n247), .ZN(n1666) );
  OAI221_X1 U1641 ( .B1(n154), .B2(n2247), .C1(n153), .C2(n2215), .A(n1074), 
        .ZN(n1067) );
  AOI22_X1 U1642 ( .A1(\REGS[29][1] ), .A2(n148), .B1(\REGS[28][1] ), .B2(n145), .ZN(n1074) );
  OAI221_X1 U1643 ( .B1(n256), .B2(n2246), .C1(n253), .C2(n2214), .A(n1684), 
        .ZN(n1677) );
  AOI22_X1 U1644 ( .A1(\REGS[29][2] ), .A2(n250), .B1(\REGS[28][2] ), .B2(n247), .ZN(n1684) );
  OAI221_X1 U1645 ( .B1(n154), .B2(n2246), .C1(n153), .C2(n2214), .A(n1092), 
        .ZN(n1085) );
  AOI22_X1 U1646 ( .A1(\REGS[29][2] ), .A2(n148), .B1(\REGS[28][2] ), .B2(n145), .ZN(n1092) );
  OAI221_X1 U1647 ( .B1(n256), .B2(n2245), .C1(n253), .C2(n2213), .A(n1702), 
        .ZN(n1695) );
  AOI22_X1 U1648 ( .A1(\REGS[29][3] ), .A2(n250), .B1(\REGS[28][3] ), .B2(n247), .ZN(n1702) );
  OAI221_X1 U1649 ( .B1(n154), .B2(n2245), .C1(n153), .C2(n2213), .A(n1110), 
        .ZN(n1103) );
  AOI22_X1 U1650 ( .A1(\REGS[29][3] ), .A2(n148), .B1(\REGS[28][3] ), .B2(n145), .ZN(n1110) );
  OAI221_X1 U1651 ( .B1(n256), .B2(n2244), .C1(n253), .C2(n2212), .A(n1720), 
        .ZN(n1713) );
  AOI22_X1 U1652 ( .A1(\REGS[29][4] ), .A2(n250), .B1(\REGS[28][4] ), .B2(n247), .ZN(n1720) );
  OAI221_X1 U1653 ( .B1(n154), .B2(n2244), .C1(n153), .C2(n2212), .A(n1128), 
        .ZN(n1121) );
  AOI22_X1 U1654 ( .A1(\REGS[29][4] ), .A2(n148), .B1(\REGS[28][4] ), .B2(n145), .ZN(n1128) );
  OAI221_X1 U1655 ( .B1(n256), .B2(n2243), .C1(n253), .C2(n2211), .A(n1738), 
        .ZN(n1731) );
  AOI22_X1 U1656 ( .A1(\REGS[29][5] ), .A2(n250), .B1(\REGS[28][5] ), .B2(n247), .ZN(n1738) );
  OAI221_X1 U1657 ( .B1(n154), .B2(n2243), .C1(n153), .C2(n2211), .A(n1146), 
        .ZN(n1139) );
  AOI22_X1 U1658 ( .A1(\REGS[29][5] ), .A2(n148), .B1(\REGS[28][5] ), .B2(n145), .ZN(n1146) );
  OAI221_X1 U1659 ( .B1(n256), .B2(n2242), .C1(n253), .C2(n2210), .A(n1756), 
        .ZN(n1749) );
  AOI22_X1 U1660 ( .A1(\REGS[29][6] ), .A2(n250), .B1(\REGS[28][6] ), .B2(n247), .ZN(n1756) );
  OAI221_X1 U1661 ( .B1(n154), .B2(n2242), .C1(n153), .C2(n2210), .A(n1164), 
        .ZN(n1157) );
  AOI22_X1 U1662 ( .A1(\REGS[29][6] ), .A2(n148), .B1(\REGS[28][6] ), .B2(n145), .ZN(n1164) );
  OAI221_X1 U1663 ( .B1(n256), .B2(n2241), .C1(n253), .C2(n2209), .A(n1774), 
        .ZN(n1767) );
  AOI22_X1 U1664 ( .A1(\REGS[29][7] ), .A2(n250), .B1(\REGS[28][7] ), .B2(n247), .ZN(n1774) );
  OAI221_X1 U1665 ( .B1(n154), .B2(n2241), .C1(n153), .C2(n2209), .A(n1182), 
        .ZN(n1175) );
  AOI22_X1 U1666 ( .A1(\REGS[29][7] ), .A2(n148), .B1(\REGS[28][7] ), .B2(n145), .ZN(n1182) );
  OAI221_X1 U1667 ( .B1(n256), .B2(n2240), .C1(n253), .C2(n2208), .A(n1792), 
        .ZN(n1785) );
  AOI22_X1 U1668 ( .A1(\REGS[29][8] ), .A2(n250), .B1(\REGS[28][8] ), .B2(n247), .ZN(n1792) );
  OAI221_X1 U1669 ( .B1(n154), .B2(n2240), .C1(n152), .C2(n2208), .A(n1200), 
        .ZN(n1193) );
  AOI22_X1 U1670 ( .A1(\REGS[29][8] ), .A2(n148), .B1(\REGS[28][8] ), .B2(n145), .ZN(n1200) );
  OAI221_X1 U1671 ( .B1(n256), .B2(n2239), .C1(n253), .C2(n2207), .A(n1810), 
        .ZN(n1803) );
  AOI22_X1 U1672 ( .A1(\REGS[29][9] ), .A2(n250), .B1(\REGS[28][9] ), .B2(n247), .ZN(n1810) );
  OAI221_X1 U1673 ( .B1(n154), .B2(n2239), .C1(n152), .C2(n2207), .A(n1218), 
        .ZN(n1211) );
  AOI22_X1 U1674 ( .A1(\REGS[29][9] ), .A2(n148), .B1(\REGS[28][9] ), .B2(n145), .ZN(n1218) );
  OAI221_X1 U1675 ( .B1(n256), .B2(n2238), .C1(n253), .C2(n2206), .A(n1837), 
        .ZN(n1821) );
  AOI22_X1 U1676 ( .A1(\REGS[29][10] ), .A2(n250), .B1(\REGS[28][10] ), .B2(
        n247), .ZN(n1837) );
  OAI221_X1 U1677 ( .B1(n154), .B2(n2238), .C1(n152), .C2(n2206), .A(n1236), 
        .ZN(n1229) );
  AOI22_X1 U1678 ( .A1(\REGS[29][10] ), .A2(n148), .B1(\REGS[28][10] ), .B2(
        n145), .ZN(n1236) );
  OAI221_X1 U1679 ( .B1(n2237), .B2(n154), .C1(n2205), .C2(n152), .A(n1254), 
        .ZN(n1247) );
  AOI22_X1 U1680 ( .A1(n148), .A2(\REGS[29][11] ), .B1(n145), .B2(
        \REGS[28][11] ), .ZN(n1254) );
  OAI221_X1 U1681 ( .B1(n2236), .B2(n155), .C1(n2204), .C2(n152), .A(n1272), 
        .ZN(n1265) );
  AOI22_X1 U1682 ( .A1(n149), .A2(\REGS[29][12] ), .B1(n146), .B2(
        \REGS[28][12] ), .ZN(n1272) );
  OAI221_X1 U1683 ( .B1(n2235), .B2(n155), .C1(n2203), .C2(n152), .A(n1290), 
        .ZN(n1283) );
  AOI22_X1 U1684 ( .A1(n149), .A2(\REGS[29][13] ), .B1(n146), .B2(
        \REGS[28][13] ), .ZN(n1290) );
  OAI221_X1 U1685 ( .B1(n2234), .B2(n155), .C1(n2202), .C2(n152), .A(n1308), 
        .ZN(n1301) );
  AOI22_X1 U1686 ( .A1(n149), .A2(\REGS[29][14] ), .B1(n146), .B2(
        \REGS[28][14] ), .ZN(n1308) );
  OAI221_X1 U1687 ( .B1(n2233), .B2(n155), .C1(n2201), .C2(n152), .A(n1326), 
        .ZN(n1319) );
  AOI22_X1 U1688 ( .A1(n149), .A2(\REGS[29][15] ), .B1(n146), .B2(
        \REGS[28][15] ), .ZN(n1326) );
  OAI221_X1 U1689 ( .B1(n2232), .B2(n155), .C1(n2200), .C2(n152), .A(n1344), 
        .ZN(n1337) );
  AOI22_X1 U1690 ( .A1(n149), .A2(\REGS[29][16] ), .B1(n146), .B2(
        \REGS[28][16] ), .ZN(n1344) );
  OAI221_X1 U1691 ( .B1(n2231), .B2(n155), .C1(n2199), .C2(n152), .A(n1362), 
        .ZN(n1355) );
  AOI22_X1 U1692 ( .A1(n149), .A2(\REGS[29][17] ), .B1(n146), .B2(
        \REGS[28][17] ), .ZN(n1362) );
  OAI221_X1 U1693 ( .B1(n2230), .B2(n155), .C1(n2198), .C2(n152), .A(n1380), 
        .ZN(n1373) );
  AOI22_X1 U1694 ( .A1(n149), .A2(\REGS[29][18] ), .B1(n146), .B2(
        \REGS[28][18] ), .ZN(n1380) );
  OAI221_X1 U1695 ( .B1(n2229), .B2(n155), .C1(n2197), .C2(n152), .A(n1398), 
        .ZN(n1391) );
  AOI22_X1 U1696 ( .A1(n149), .A2(\REGS[29][19] ), .B1(n146), .B2(
        \REGS[28][19] ), .ZN(n1398) );
  OAI221_X1 U1697 ( .B1(n257), .B2(n2229), .C1(n254), .C2(n2197), .A(n744), 
        .ZN(n737) );
  AOI22_X1 U1698 ( .A1(\REGS[29][19] ), .A2(n251), .B1(\REGS[28][19] ), .B2(
        n248), .ZN(n744) );
  OAI221_X1 U1699 ( .B1(n2228), .B2(n155), .C1(n2196), .C2(n151), .A(n1416), 
        .ZN(n1409) );
  AOI22_X1 U1700 ( .A1(n149), .A2(\REGS[29][20] ), .B1(n146), .B2(
        \REGS[28][20] ), .ZN(n1416) );
  OAI221_X1 U1701 ( .B1(n257), .B2(n2228), .C1(n254), .C2(n2196), .A(n762), 
        .ZN(n755) );
  AOI22_X1 U1702 ( .A1(\REGS[29][20] ), .A2(n251), .B1(\REGS[28][20] ), .B2(
        n248), .ZN(n762) );
  OAI221_X1 U1703 ( .B1(n2227), .B2(n155), .C1(n2195), .C2(n151), .A(n1434), 
        .ZN(n1427) );
  AOI22_X1 U1704 ( .A1(n149), .A2(\REGS[29][21] ), .B1(n146), .B2(
        \REGS[28][21] ), .ZN(n1434) );
  OAI221_X1 U1705 ( .B1(n257), .B2(n2227), .C1(n254), .C2(n2195), .A(n780), 
        .ZN(n773) );
  AOI22_X1 U1706 ( .A1(\REGS[29][21] ), .A2(n251), .B1(\REGS[28][21] ), .B2(
        n248), .ZN(n780) );
  OAI221_X1 U1707 ( .B1(n2226), .B2(n155), .C1(n2194), .C2(n151), .A(n1452), 
        .ZN(n1445) );
  AOI22_X1 U1708 ( .A1(n149), .A2(\REGS[29][22] ), .B1(n146), .B2(
        \REGS[28][22] ), .ZN(n1452) );
  OAI221_X1 U1709 ( .B1(n257), .B2(n2226), .C1(n254), .C2(n2194), .A(n798), 
        .ZN(n791) );
  AOI22_X1 U1710 ( .A1(\REGS[29][22] ), .A2(n251), .B1(\REGS[28][22] ), .B2(
        n248), .ZN(n798) );
  OAI221_X1 U1711 ( .B1(n2225), .B2(n155), .C1(n2193), .C2(n151), .A(n1470), 
        .ZN(n1463) );
  AOI22_X1 U1712 ( .A1(n149), .A2(\REGS[29][23] ), .B1(n146), .B2(
        \REGS[28][23] ), .ZN(n1470) );
  OAI221_X1 U1713 ( .B1(n257), .B2(n2225), .C1(n254), .C2(n2193), .A(n816), 
        .ZN(n809) );
  AOI22_X1 U1714 ( .A1(\REGS[29][23] ), .A2(n251), .B1(\REGS[28][23] ), .B2(
        n248), .ZN(n816) );
  OAI221_X1 U1715 ( .B1(n2224), .B2(n155), .C1(n2192), .C2(n151), .A(n1488), 
        .ZN(n1481) );
  AOI22_X1 U1716 ( .A1(n149), .A2(\REGS[29][24] ), .B1(n146), .B2(
        \REGS[28][24] ), .ZN(n1488) );
  OAI221_X1 U1717 ( .B1(n257), .B2(n2224), .C1(n254), .C2(n2192), .A(n834), 
        .ZN(n827) );
  AOI22_X1 U1718 ( .A1(\REGS[29][24] ), .A2(n251), .B1(\REGS[28][24] ), .B2(
        n248), .ZN(n834) );
  OAI221_X1 U1719 ( .B1(n257), .B2(n2223), .C1(n254), .C2(n2191), .A(n852), 
        .ZN(n845) );
  AOI22_X1 U1720 ( .A1(\REGS[29][25] ), .A2(n251), .B1(\REGS[28][25] ), .B2(
        n248), .ZN(n852) );
  OAI221_X1 U1721 ( .B1(n257), .B2(n2222), .C1(n254), .C2(n2190), .A(n870), 
        .ZN(n863) );
  AOI22_X1 U1722 ( .A1(\REGS[29][26] ), .A2(n251), .B1(\REGS[28][26] ), .B2(
        n248), .ZN(n870) );
  OAI221_X1 U1723 ( .B1(n257), .B2(n2221), .C1(n254), .C2(n2189), .A(n888), 
        .ZN(n881) );
  AOI22_X1 U1724 ( .A1(\REGS[29][27] ), .A2(n251), .B1(\REGS[28][27] ), .B2(
        n248), .ZN(n888) );
  OAI221_X1 U1725 ( .B1(n257), .B2(n2220), .C1(n254), .C2(n2188), .A(n906), 
        .ZN(n899) );
  AOI22_X1 U1726 ( .A1(\REGS[29][28] ), .A2(n251), .B1(\REGS[28][28] ), .B2(
        n248), .ZN(n906) );
  OAI221_X1 U1727 ( .B1(n257), .B2(n2219), .C1(n254), .C2(n2187), .A(n924), 
        .ZN(n917) );
  AOI22_X1 U1728 ( .A1(\REGS[29][29] ), .A2(n251), .B1(\REGS[28][29] ), .B2(
        n248), .ZN(n924) );
  OAI221_X1 U1729 ( .B1(n257), .B2(n2218), .C1(n254), .C2(n2186), .A(n942), 
        .ZN(n935) );
  AOI22_X1 U1730 ( .A1(\REGS[29][30] ), .A2(n251), .B1(\REGS[28][30] ), .B2(
        n248), .ZN(n942) );
  OAI221_X1 U1731 ( .B1(n256), .B2(n2217), .C1(n253), .C2(n2185), .A(n960), 
        .ZN(n953) );
  AOI22_X1 U1732 ( .A1(\REGS[29][31] ), .A2(n250), .B1(\REGS[28][31] ), .B2(
        n247), .ZN(n960) );
  AOI21_X1 U1733 ( .B1(n198), .B2(WE), .A(n391), .ZN(n1002) );
  AOI22_X1 U1734 ( .A1(\REGS[15][11] ), .A2(n204), .B1(\REGS[14][11] ), .B2(
        n201), .ZN(n606) );
  AOI22_X1 U1735 ( .A1(\REGS[15][12] ), .A2(n204), .B1(\REGS[14][12] ), .B2(
        n201), .ZN(n626) );
  AOI22_X1 U1736 ( .A1(\REGS[15][13] ), .A2(n204), .B1(\REGS[14][13] ), .B2(
        n201), .ZN(n644) );
  AOI22_X1 U1737 ( .A1(\REGS[15][14] ), .A2(n204), .B1(\REGS[14][14] ), .B2(
        n201), .ZN(n662) );
  AOI22_X1 U1738 ( .A1(\REGS[15][15] ), .A2(n204), .B1(\REGS[14][15] ), .B2(
        n201), .ZN(n680) );
  AOI22_X1 U1739 ( .A1(\REGS[15][16] ), .A2(n204), .B1(\REGS[14][16] ), .B2(
        n201), .ZN(n698) );
  AOI22_X1 U1740 ( .A1(\REGS[15][17] ), .A2(n204), .B1(\REGS[14][17] ), .B2(
        n201), .ZN(n716) );
  AOI22_X1 U1741 ( .A1(\REGS[15][18] ), .A2(n204), .B1(\REGS[14][18] ), .B2(
        n201), .ZN(n734) );
  AOI22_X1 U1742 ( .A1(\REGS[15][0] ), .A2(n202), .B1(\REGS[14][0] ), .B2(n199), .ZN(n1656) );
  AOI22_X1 U1743 ( .A1(\REGS[15][0] ), .A2(n100), .B1(\REGS[14][0] ), .B2(n97), 
        .ZN(n1062) );
  AOI22_X1 U1744 ( .A1(\REGS[15][1] ), .A2(n202), .B1(\REGS[14][1] ), .B2(n199), .ZN(n1674) );
  AOI22_X1 U1745 ( .A1(\REGS[15][1] ), .A2(n100), .B1(\REGS[14][1] ), .B2(n97), 
        .ZN(n1082) );
  AOI22_X1 U1746 ( .A1(\REGS[15][2] ), .A2(n202), .B1(\REGS[14][2] ), .B2(n199), .ZN(n1692) );
  AOI22_X1 U1747 ( .A1(\REGS[15][2] ), .A2(n100), .B1(\REGS[14][2] ), .B2(n97), 
        .ZN(n1100) );
  AOI22_X1 U1748 ( .A1(\REGS[15][3] ), .A2(n202), .B1(\REGS[14][3] ), .B2(n199), .ZN(n1710) );
  AOI22_X1 U1749 ( .A1(\REGS[15][3] ), .A2(n100), .B1(\REGS[14][3] ), .B2(n97), 
        .ZN(n1118) );
  AOI22_X1 U1750 ( .A1(\REGS[15][4] ), .A2(n202), .B1(\REGS[14][4] ), .B2(n199), .ZN(n1728) );
  AOI22_X1 U1751 ( .A1(\REGS[15][4] ), .A2(n100), .B1(\REGS[14][4] ), .B2(n97), 
        .ZN(n1136) );
  AOI22_X1 U1752 ( .A1(\REGS[15][5] ), .A2(n202), .B1(\REGS[14][5] ), .B2(n199), .ZN(n1746) );
  AOI22_X1 U1753 ( .A1(\REGS[15][5] ), .A2(n100), .B1(\REGS[14][5] ), .B2(n97), 
        .ZN(n1154) );
  AOI22_X1 U1754 ( .A1(\REGS[15][6] ), .A2(n202), .B1(\REGS[14][6] ), .B2(n199), .ZN(n1764) );
  AOI22_X1 U1755 ( .A1(\REGS[15][6] ), .A2(n100), .B1(\REGS[14][6] ), .B2(n97), 
        .ZN(n1172) );
  AOI22_X1 U1756 ( .A1(\REGS[15][7] ), .A2(n202), .B1(\REGS[14][7] ), .B2(n199), .ZN(n1782) );
  AOI22_X1 U1757 ( .A1(\REGS[15][7] ), .A2(n100), .B1(\REGS[14][7] ), .B2(n97), 
        .ZN(n1190) );
  AOI22_X1 U1758 ( .A1(\REGS[15][8] ), .A2(n202), .B1(\REGS[14][8] ), .B2(n199), .ZN(n1800) );
  AOI22_X1 U1759 ( .A1(\REGS[15][8] ), .A2(n100), .B1(\REGS[14][8] ), .B2(n97), 
        .ZN(n1208) );
  AOI22_X1 U1760 ( .A1(\REGS[15][9] ), .A2(n202), .B1(\REGS[14][9] ), .B2(n199), .ZN(n1818) );
  AOI22_X1 U1761 ( .A1(\REGS[15][9] ), .A2(n100), .B1(\REGS[14][9] ), .B2(n97), 
        .ZN(n1226) );
  AOI22_X1 U1762 ( .A1(\REGS[15][10] ), .A2(n202), .B1(\REGS[14][10] ), .B2(
        n199), .ZN(n1851) );
  AOI22_X1 U1763 ( .A1(\REGS[15][10] ), .A2(n100), .B1(\REGS[14][10] ), .B2(
        n97), .ZN(n1244) );
  AOI22_X1 U1764 ( .A1(n100), .A2(\REGS[15][11] ), .B1(n97), .B2(
        \REGS[14][11] ), .ZN(n1262) );
  AOI22_X1 U1765 ( .A1(n101), .A2(\REGS[15][12] ), .B1(n98), .B2(
        \REGS[14][12] ), .ZN(n1280) );
  AOI22_X1 U1766 ( .A1(n101), .A2(\REGS[15][13] ), .B1(n98), .B2(
        \REGS[14][13] ), .ZN(n1298) );
  AOI22_X1 U1767 ( .A1(n101), .A2(\REGS[15][14] ), .B1(n98), .B2(
        \REGS[14][14] ), .ZN(n1316) );
  AOI22_X1 U1768 ( .A1(n101), .A2(\REGS[15][15] ), .B1(n98), .B2(
        \REGS[14][15] ), .ZN(n1334) );
  AOI22_X1 U1769 ( .A1(n101), .A2(\REGS[15][16] ), .B1(n98), .B2(
        \REGS[14][16] ), .ZN(n1352) );
  AOI22_X1 U1770 ( .A1(n101), .A2(\REGS[15][17] ), .B1(n98), .B2(
        \REGS[14][17] ), .ZN(n1370) );
  AOI22_X1 U1771 ( .A1(n101), .A2(\REGS[15][18] ), .B1(n98), .B2(
        \REGS[14][18] ), .ZN(n1388) );
  AOI22_X1 U1772 ( .A1(n101), .A2(\REGS[15][19] ), .B1(n98), .B2(
        \REGS[14][19] ), .ZN(n1406) );
  AOI22_X1 U1773 ( .A1(\REGS[15][19] ), .A2(n203), .B1(\REGS[14][19] ), .B2(
        n200), .ZN(n752) );
  AOI22_X1 U1774 ( .A1(n101), .A2(\REGS[15][20] ), .B1(n98), .B2(
        \REGS[14][20] ), .ZN(n1424) );
  AOI22_X1 U1775 ( .A1(\REGS[15][20] ), .A2(n203), .B1(\REGS[14][20] ), .B2(
        n200), .ZN(n770) );
  AOI22_X1 U1776 ( .A1(n101), .A2(\REGS[15][21] ), .B1(n98), .B2(
        \REGS[14][21] ), .ZN(n1442) );
  AOI22_X1 U1777 ( .A1(\REGS[15][21] ), .A2(n203), .B1(\REGS[14][21] ), .B2(
        n200), .ZN(n788) );
  AOI22_X1 U1778 ( .A1(n101), .A2(\REGS[15][22] ), .B1(n98), .B2(
        \REGS[14][22] ), .ZN(n1460) );
  AOI22_X1 U1779 ( .A1(\REGS[15][22] ), .A2(n203), .B1(\REGS[14][22] ), .B2(
        n200), .ZN(n806) );
  AOI22_X1 U1780 ( .A1(n101), .A2(\REGS[15][23] ), .B1(n98), .B2(
        \REGS[14][23] ), .ZN(n1478) );
  AOI22_X1 U1781 ( .A1(\REGS[15][23] ), .A2(n203), .B1(\REGS[14][23] ), .B2(
        n200), .ZN(n824) );
  AOI22_X1 U1782 ( .A1(n101), .A2(\REGS[15][24] ), .B1(n98), .B2(
        \REGS[14][24] ), .ZN(n1496) );
  AOI22_X1 U1783 ( .A1(\REGS[15][24] ), .A2(n203), .B1(\REGS[14][24] ), .B2(
        n200), .ZN(n842) );
  AOI22_X1 U1784 ( .A1(n102), .A2(\REGS[15][25] ), .B1(n99), .B2(
        \REGS[14][25] ), .ZN(n1514) );
  AOI22_X1 U1785 ( .A1(\REGS[15][25] ), .A2(n203), .B1(\REGS[14][25] ), .B2(
        n200), .ZN(n860) );
  AOI22_X1 U1786 ( .A1(n102), .A2(\REGS[15][26] ), .B1(n99), .B2(
        \REGS[14][26] ), .ZN(n1532) );
  AOI22_X1 U1787 ( .A1(\REGS[15][26] ), .A2(n203), .B1(\REGS[14][26] ), .B2(
        n200), .ZN(n878) );
  AOI22_X1 U1788 ( .A1(n102), .A2(\REGS[15][27] ), .B1(n99), .B2(
        \REGS[14][27] ), .ZN(n1550) );
  AOI22_X1 U1789 ( .A1(\REGS[15][27] ), .A2(n203), .B1(\REGS[14][27] ), .B2(
        n200), .ZN(n896) );
  AOI22_X1 U1790 ( .A1(n102), .A2(\REGS[15][28] ), .B1(n99), .B2(
        \REGS[14][28] ), .ZN(n1568) );
  AOI22_X1 U1791 ( .A1(\REGS[15][28] ), .A2(n203), .B1(\REGS[14][28] ), .B2(
        n200), .ZN(n914) );
  AOI22_X1 U1792 ( .A1(n102), .A2(\REGS[15][29] ), .B1(n99), .B2(
        \REGS[14][29] ), .ZN(n1586) );
  AOI22_X1 U1793 ( .A1(\REGS[15][29] ), .A2(n203), .B1(\REGS[14][29] ), .B2(
        n200), .ZN(n932) );
  AOI22_X1 U1794 ( .A1(n102), .A2(\REGS[15][30] ), .B1(n99), .B2(
        \REGS[14][30] ), .ZN(n1604) );
  AOI22_X1 U1795 ( .A1(\REGS[15][30] ), .A2(n203), .B1(\REGS[14][30] ), .B2(
        n200), .ZN(n950) );
  AOI22_X1 U1796 ( .A1(n102), .A2(\REGS[15][31] ), .B1(n99), .B2(
        \REGS[14][31] ), .ZN(n1637) );
  AOI22_X1 U1797 ( .A1(\REGS[15][31] ), .A2(n202), .B1(\REGS[14][31] ), .B2(
        n199), .ZN(n968) );
  NAND2_X1 U1798 ( .A1(DATA_IN[20]), .A2(n389), .ZN(n981) );
  NAND2_X1 U1799 ( .A1(DATA_IN[21]), .A2(n388), .ZN(n980) );
  NAND2_X1 U1800 ( .A1(DATA_IN[22]), .A2(n389), .ZN(n979) );
  NAND2_X1 U1801 ( .A1(DATA_IN[23]), .A2(n390), .ZN(n978) );
  NAND2_X1 U1802 ( .A1(DATA_IN[24]), .A2(n389), .ZN(n977) );
  NAND2_X1 U1803 ( .A1(DATA_IN[25]), .A2(n388), .ZN(n976) );
  NAND2_X1 U1804 ( .A1(DATA_IN[26]), .A2(n389), .ZN(n975) );
  NAND2_X1 U1805 ( .A1(DATA_IN[27]), .A2(n390), .ZN(n974) );
  NAND2_X1 U1806 ( .A1(DATA_IN[28]), .A2(n390), .ZN(n973) );
  NAND2_X1 U1807 ( .A1(DATA_IN[29]), .A2(n388), .ZN(n972) );
  NAND2_X1 U1808 ( .A1(DATA_IN[30]), .A2(n389), .ZN(n971) );
  NAND2_X1 U1809 ( .A1(DATA_IN[31]), .A2(n390), .ZN(n970) );
  AND2_X1 U1810 ( .A1(ADDR_RD2[0]), .A2(n1624), .ZN(n1622) );
  AND2_X1 U1811 ( .A1(ADDR_RD1[0]), .A2(n1838), .ZN(n1836) );
  NOR2_X1 U1812 ( .A1(ADDR_RD2[3]), .A2(ADDR_RD2[4]), .ZN(n1633) );
  NOR2_X1 U1813 ( .A1(n407), .A2(ADDR_RD2[4]), .ZN(n1638) );
  NOR2_X1 U1814 ( .A1(ADDR_RD1[3]), .A2(ADDR_RD1[4]), .ZN(n1847) );
  NOR2_X1 U1815 ( .A1(n403), .A2(ADDR_RD1[4]), .ZN(n1852) );
  AND2_X1 U1816 ( .A1(n1619), .A2(ADDR_RD2[0]), .ZN(n1614) );
  AND2_X1 U1817 ( .A1(n1633), .A2(ADDR_RD2[0]), .ZN(n1631) );
  AND2_X1 U1818 ( .A1(n1638), .A2(ADDR_RD2[0]), .ZN(n1636) );
  AND2_X1 U1819 ( .A1(n1833), .A2(ADDR_RD1[0]), .ZN(n1828) );
  AND2_X1 U1820 ( .A1(n1847), .A2(ADDR_RD1[0]), .ZN(n1845) );
  AND2_X1 U1821 ( .A1(n1852), .A2(ADDR_RD1[0]), .ZN(n1850) );
  NAND2_X1 U1822 ( .A1(DATA_IN[8]), .A2(n388), .ZN(n993) );
  NAND2_X1 U1823 ( .A1(DATA_IN[9]), .A2(n388), .ZN(n992) );
  NAND2_X1 U1824 ( .A1(DATA_IN[10]), .A2(n388), .ZN(n991) );
  NAND2_X1 U1825 ( .A1(DATA_IN[11]), .A2(n388), .ZN(n990) );
  NAND2_X1 U1826 ( .A1(DATA_IN[12]), .A2(n388), .ZN(n989) );
  NAND2_X1 U1827 ( .A1(DATA_IN[13]), .A2(n388), .ZN(n988) );
  NAND2_X1 U1828 ( .A1(DATA_IN[14]), .A2(n388), .ZN(n987) );
  NAND2_X1 U1829 ( .A1(DATA_IN[15]), .A2(n388), .ZN(n986) );
  NAND2_X1 U1830 ( .A1(DATA_IN[16]), .A2(n388), .ZN(n985) );
  NAND2_X1 U1831 ( .A1(DATA_IN[17]), .A2(n388), .ZN(n984) );
  NAND2_X1 U1832 ( .A1(DATA_IN[18]), .A2(n388), .ZN(n983) );
  NAND2_X1 U1833 ( .A1(DATA_IN[19]), .A2(n388), .ZN(n982) );
  NAND2_X1 U1834 ( .A1(DATA_IN[0]), .A2(n389), .ZN(n1001) );
  NAND2_X1 U1835 ( .A1(DATA_IN[1]), .A2(n389), .ZN(n1000) );
  NAND2_X1 U1836 ( .A1(DATA_IN[2]), .A2(n389), .ZN(n999) );
  NAND2_X1 U1837 ( .A1(DATA_IN[3]), .A2(n389), .ZN(n998) );
  NAND2_X1 U1838 ( .A1(DATA_IN[4]), .A2(n389), .ZN(n997) );
  NAND2_X1 U1839 ( .A1(DATA_IN[5]), .A2(n389), .ZN(n996) );
  NAND2_X1 U1840 ( .A1(DATA_IN[6]), .A2(n389), .ZN(n995) );
  NAND2_X1 U1841 ( .A1(DATA_IN[7]), .A2(n389), .ZN(n994) );
  INV_X1 U1842 ( .A(ADDR_RD2[0]), .ZN(n410) );
  INV_X1 U1843 ( .A(ADDR_RD1[0]), .ZN(n406) );
  INV_X1 U1844 ( .A(ADDR_RD2[1]), .ZN(n409) );
  INV_X1 U1845 ( .A(ADDR_RD2[2]), .ZN(n408) );
  INV_X1 U1846 ( .A(ADDR_RD1[1]), .ZN(n405) );
  INV_X1 U1847 ( .A(ADDR_RD1[2]), .ZN(n404) );
  INV_X1 U1848 ( .A(\REGS[17][11] ), .ZN(n2045) );
  INV_X1 U1849 ( .A(\REGS[21][11] ), .ZN(n2109) );
  INV_X1 U1850 ( .A(\REGS[25][11] ), .ZN(n2173) );
  INV_X1 U1851 ( .A(\REGS[31][11] ), .ZN(n2237) );
  INV_X1 U1852 ( .A(\REGS[1][11] ), .ZN(n495) );
  INV_X1 U1853 ( .A(\REGS[5][11] ), .ZN(n1853) );
  INV_X1 U1854 ( .A(\REGS[9][11] ), .ZN(n1917) );
  INV_X1 U1855 ( .A(\REGS[13][11] ), .ZN(n1981) );
  INV_X1 U1856 ( .A(\REGS[17][12] ), .ZN(n2044) );
  INV_X1 U1857 ( .A(\REGS[21][12] ), .ZN(n2108) );
  INV_X1 U1858 ( .A(\REGS[25][12] ), .ZN(n2172) );
  INV_X1 U1859 ( .A(\REGS[31][12] ), .ZN(n2236) );
  INV_X1 U1860 ( .A(\REGS[1][12] ), .ZN(n494) );
  INV_X1 U1861 ( .A(\REGS[5][12] ), .ZN(n558) );
  INV_X1 U1862 ( .A(\REGS[9][12] ), .ZN(n1916) );
  INV_X1 U1863 ( .A(\REGS[13][12] ), .ZN(n1980) );
  INV_X1 U1864 ( .A(\REGS[17][13] ), .ZN(n2043) );
  INV_X1 U1865 ( .A(\REGS[21][13] ), .ZN(n2107) );
  INV_X1 U1866 ( .A(\REGS[25][13] ), .ZN(n2171) );
  INV_X1 U1867 ( .A(\REGS[31][13] ), .ZN(n2235) );
  INV_X1 U1868 ( .A(\REGS[1][13] ), .ZN(n493) );
  INV_X1 U1869 ( .A(\REGS[5][13] ), .ZN(n557) );
  INV_X1 U1870 ( .A(\REGS[9][13] ), .ZN(n1915) );
  INV_X1 U1871 ( .A(\REGS[13][13] ), .ZN(n1979) );
  INV_X1 U1872 ( .A(\REGS[17][14] ), .ZN(n2042) );
  INV_X1 U1873 ( .A(\REGS[21][14] ), .ZN(n2106) );
  INV_X1 U1874 ( .A(\REGS[25][14] ), .ZN(n2170) );
  INV_X1 U1875 ( .A(\REGS[31][14] ), .ZN(n2234) );
  INV_X1 U1876 ( .A(\REGS[1][14] ), .ZN(n492) );
  INV_X1 U1877 ( .A(\REGS[5][14] ), .ZN(n556) );
  INV_X1 U1878 ( .A(\REGS[9][14] ), .ZN(n1914) );
  INV_X1 U1879 ( .A(\REGS[13][14] ), .ZN(n1978) );
  INV_X1 U1880 ( .A(\REGS[17][15] ), .ZN(n2041) );
  INV_X1 U1881 ( .A(\REGS[21][15] ), .ZN(n2105) );
  INV_X1 U1882 ( .A(\REGS[25][15] ), .ZN(n2169) );
  INV_X1 U1883 ( .A(\REGS[31][15] ), .ZN(n2233) );
  INV_X1 U1884 ( .A(\REGS[1][15] ), .ZN(n491) );
  INV_X1 U1885 ( .A(\REGS[5][15] ), .ZN(n555) );
  INV_X1 U1886 ( .A(\REGS[9][15] ), .ZN(n1913) );
  INV_X1 U1887 ( .A(\REGS[13][15] ), .ZN(n1977) );
  INV_X1 U1888 ( .A(\REGS[17][16] ), .ZN(n2040) );
  INV_X1 U1889 ( .A(\REGS[21][16] ), .ZN(n2104) );
  INV_X1 U1890 ( .A(\REGS[25][16] ), .ZN(n2168) );
  INV_X1 U1891 ( .A(\REGS[31][16] ), .ZN(n2232) );
  INV_X1 U1892 ( .A(\REGS[1][16] ), .ZN(n490) );
  INV_X1 U1893 ( .A(\REGS[5][16] ), .ZN(n554) );
  INV_X1 U1894 ( .A(\REGS[9][16] ), .ZN(n1912) );
  INV_X1 U1895 ( .A(\REGS[13][16] ), .ZN(n1976) );
  INV_X1 U1896 ( .A(\REGS[17][17] ), .ZN(n2039) );
  INV_X1 U1897 ( .A(\REGS[21][17] ), .ZN(n2103) );
  INV_X1 U1898 ( .A(\REGS[25][17] ), .ZN(n2167) );
  INV_X1 U1899 ( .A(\REGS[31][17] ), .ZN(n2231) );
  INV_X1 U1900 ( .A(\REGS[1][17] ), .ZN(n489) );
  INV_X1 U1901 ( .A(\REGS[5][17] ), .ZN(n553) );
  INV_X1 U1902 ( .A(\REGS[9][17] ), .ZN(n1911) );
  INV_X1 U1903 ( .A(\REGS[13][17] ), .ZN(n1975) );
  INV_X1 U1904 ( .A(\REGS[17][18] ), .ZN(n2038) );
  INV_X1 U1905 ( .A(\REGS[21][18] ), .ZN(n2102) );
  INV_X1 U1906 ( .A(\REGS[25][18] ), .ZN(n2166) );
  INV_X1 U1907 ( .A(\REGS[31][18] ), .ZN(n2230) );
  INV_X1 U1908 ( .A(\REGS[1][18] ), .ZN(n488) );
  INV_X1 U1909 ( .A(\REGS[5][18] ), .ZN(n552) );
  INV_X1 U1910 ( .A(\REGS[9][18] ), .ZN(n1910) );
  INV_X1 U1911 ( .A(\REGS[13][18] ), .ZN(n1974) );
  INV_X1 U1912 ( .A(\REGS[17][19] ), .ZN(n2037) );
  INV_X1 U1913 ( .A(\REGS[21][19] ), .ZN(n2101) );
  INV_X1 U1914 ( .A(\REGS[25][19] ), .ZN(n2165) );
  INV_X1 U1915 ( .A(\REGS[31][19] ), .ZN(n2229) );
  INV_X1 U1916 ( .A(\REGS[1][19] ), .ZN(n487) );
  INV_X1 U1917 ( .A(\REGS[5][19] ), .ZN(n551) );
  INV_X1 U1918 ( .A(\REGS[9][19] ), .ZN(n1909) );
  INV_X1 U1919 ( .A(\REGS[13][19] ), .ZN(n1973) );
  INV_X1 U1920 ( .A(\REGS[17][20] ), .ZN(n2036) );
  INV_X1 U1921 ( .A(\REGS[21][20] ), .ZN(n2100) );
  INV_X1 U1922 ( .A(\REGS[25][20] ), .ZN(n2164) );
  INV_X1 U1923 ( .A(\REGS[31][20] ), .ZN(n2228) );
  INV_X1 U1924 ( .A(\REGS[1][20] ), .ZN(n486) );
  INV_X1 U1925 ( .A(\REGS[5][20] ), .ZN(n550) );
  INV_X1 U1926 ( .A(\REGS[9][20] ), .ZN(n1908) );
  INV_X1 U1927 ( .A(\REGS[13][20] ), .ZN(n1972) );
  INV_X1 U1928 ( .A(\REGS[17][21] ), .ZN(n2035) );
  INV_X1 U1929 ( .A(\REGS[21][21] ), .ZN(n2099) );
  INV_X1 U1930 ( .A(\REGS[25][21] ), .ZN(n2163) );
  INV_X1 U1931 ( .A(\REGS[31][21] ), .ZN(n2227) );
  INV_X1 U1932 ( .A(\REGS[1][21] ), .ZN(n485) );
  INV_X1 U1933 ( .A(\REGS[5][21] ), .ZN(n549) );
  INV_X1 U1934 ( .A(\REGS[9][21] ), .ZN(n1907) );
  INV_X1 U1935 ( .A(\REGS[13][21] ), .ZN(n1971) );
  INV_X1 U1936 ( .A(\REGS[17][22] ), .ZN(n2034) );
  INV_X1 U1937 ( .A(\REGS[21][22] ), .ZN(n2098) );
  INV_X1 U1938 ( .A(\REGS[25][22] ), .ZN(n2162) );
  INV_X1 U1939 ( .A(\REGS[31][22] ), .ZN(n2226) );
  INV_X1 U1940 ( .A(\REGS[1][22] ), .ZN(n484) );
  INV_X1 U1941 ( .A(\REGS[5][22] ), .ZN(n548) );
  INV_X1 U1942 ( .A(\REGS[9][22] ), .ZN(n1906) );
  INV_X1 U1943 ( .A(\REGS[13][22] ), .ZN(n1970) );
  INV_X1 U1944 ( .A(\REGS[17][23] ), .ZN(n2033) );
  INV_X1 U1945 ( .A(\REGS[21][23] ), .ZN(n2097) );
  INV_X1 U1946 ( .A(\REGS[25][23] ), .ZN(n2161) );
  INV_X1 U1947 ( .A(\REGS[31][23] ), .ZN(n2225) );
  INV_X1 U1948 ( .A(\REGS[1][23] ), .ZN(n483) );
  INV_X1 U1949 ( .A(\REGS[5][23] ), .ZN(n547) );
  INV_X1 U1950 ( .A(\REGS[9][23] ), .ZN(n1905) );
  INV_X1 U1951 ( .A(\REGS[13][23] ), .ZN(n1969) );
  INV_X1 U1952 ( .A(\REGS[17][24] ), .ZN(n2032) );
  INV_X1 U1953 ( .A(\REGS[21][24] ), .ZN(n2096) );
  INV_X1 U1954 ( .A(\REGS[25][24] ), .ZN(n2160) );
  INV_X1 U1955 ( .A(\REGS[31][24] ), .ZN(n2224) );
  INV_X1 U1956 ( .A(\REGS[1][24] ), .ZN(n482) );
  INV_X1 U1957 ( .A(\REGS[5][24] ), .ZN(n546) );
  INV_X1 U1958 ( .A(\REGS[9][24] ), .ZN(n1904) );
  INV_X1 U1959 ( .A(\REGS[13][24] ), .ZN(n1968) );
  INV_X1 U1960 ( .A(\REGS[17][25] ), .ZN(n2031) );
  INV_X1 U1961 ( .A(\REGS[21][25] ), .ZN(n2095) );
  INV_X1 U1962 ( .A(\REGS[25][25] ), .ZN(n2159) );
  INV_X1 U1963 ( .A(\REGS[31][25] ), .ZN(n2223) );
  INV_X1 U1964 ( .A(\REGS[1][25] ), .ZN(n481) );
  INV_X1 U1965 ( .A(\REGS[5][25] ), .ZN(n545) );
  INV_X1 U1966 ( .A(\REGS[9][25] ), .ZN(n1903) );
  INV_X1 U1967 ( .A(\REGS[13][25] ), .ZN(n1967) );
  INV_X1 U1968 ( .A(\REGS[17][26] ), .ZN(n2030) );
  INV_X1 U1969 ( .A(\REGS[21][26] ), .ZN(n2094) );
  INV_X1 U1982 ( .A(\REGS[25][26] ), .ZN(n2158) );
  INV_X1 U1983 ( .A(\REGS[31][26] ), .ZN(n2222) );
  INV_X1 U1984 ( .A(\REGS[1][26] ), .ZN(n480) );
  INV_X1 U1985 ( .A(\REGS[5][26] ), .ZN(n544) );
  INV_X1 U1986 ( .A(\REGS[9][26] ), .ZN(n1902) );
  INV_X1 U1987 ( .A(\REGS[13][26] ), .ZN(n1966) );
  INV_X1 U1988 ( .A(\REGS[17][27] ), .ZN(n2029) );
  INV_X1 U1989 ( .A(\REGS[21][27] ), .ZN(n2093) );
  INV_X1 U1990 ( .A(\REGS[25][27] ), .ZN(n2157) );
  INV_X1 U1991 ( .A(\REGS[31][27] ), .ZN(n2221) );
  INV_X1 U1992 ( .A(\REGS[1][27] ), .ZN(n479) );
  INV_X1 U1993 ( .A(\REGS[5][27] ), .ZN(n543) );
  INV_X1 U1994 ( .A(\REGS[9][27] ), .ZN(n1901) );
  INV_X1 U1995 ( .A(\REGS[13][27] ), .ZN(n1965) );
  INV_X1 U1996 ( .A(\REGS[17][28] ), .ZN(n2028) );
  INV_X1 U1997 ( .A(\REGS[21][28] ), .ZN(n2092) );
  INV_X1 U1998 ( .A(\REGS[25][28] ), .ZN(n2156) );
  INV_X1 U1999 ( .A(\REGS[31][28] ), .ZN(n2220) );
  INV_X1 U2000 ( .A(\REGS[1][28] ), .ZN(n478) );
  INV_X1 U2001 ( .A(\REGS[5][28] ), .ZN(n542) );
  INV_X1 U2002 ( .A(\REGS[9][28] ), .ZN(n1900) );
  INV_X1 U2003 ( .A(\REGS[13][28] ), .ZN(n1964) );
  INV_X1 U2004 ( .A(\REGS[17][29] ), .ZN(n2027) );
  INV_X1 U2005 ( .A(\REGS[21][29] ), .ZN(n2091) );
  INV_X1 U2006 ( .A(\REGS[25][29] ), .ZN(n2155) );
  INV_X1 U2007 ( .A(\REGS[31][29] ), .ZN(n2219) );
  INV_X1 U2008 ( .A(\REGS[1][29] ), .ZN(n477) );
  INV_X1 U2009 ( .A(\REGS[5][29] ), .ZN(n541) );
  INV_X1 U2010 ( .A(\REGS[9][29] ), .ZN(n1899) );
  INV_X1 U2011 ( .A(\REGS[13][29] ), .ZN(n1963) );
  INV_X1 U2012 ( .A(\REGS[17][30] ), .ZN(n2026) );
  INV_X1 U2013 ( .A(\REGS[21][30] ), .ZN(n2090) );
  INV_X1 U2014 ( .A(\REGS[25][30] ), .ZN(n2154) );
  INV_X1 U2015 ( .A(\REGS[31][30] ), .ZN(n2218) );
  INV_X1 U2016 ( .A(\REGS[1][30] ), .ZN(n476) );
  INV_X1 U2017 ( .A(\REGS[5][30] ), .ZN(n540) );
  INV_X1 U2018 ( .A(\REGS[9][30] ), .ZN(n1898) );
  INV_X1 U2019 ( .A(\REGS[13][30] ), .ZN(n1962) );
  INV_X1 U2020 ( .A(\REGS[17][31] ), .ZN(n2025) );
  INV_X1 U2021 ( .A(\REGS[21][31] ), .ZN(n2089) );
  INV_X1 U2022 ( .A(\REGS[25][31] ), .ZN(n2153) );
  INV_X1 U2023 ( .A(\REGS[31][31] ), .ZN(n2217) );
  INV_X1 U2024 ( .A(\REGS[1][31] ), .ZN(n475) );
  INV_X1 U2025 ( .A(\REGS[5][31] ), .ZN(n539) );
  INV_X1 U2026 ( .A(\REGS[9][31] ), .ZN(n1897) );
  INV_X1 U2027 ( .A(\REGS[13][31] ), .ZN(n1961) );
  INV_X1 U2028 ( .A(\REGS[16][0] ), .ZN(n2024) );
  INV_X1 U2029 ( .A(\REGS[20][0] ), .ZN(n2088) );
  INV_X1 U2030 ( .A(\REGS[24][0] ), .ZN(n2152) );
  INV_X1 U2031 ( .A(\REGS[30][0] ), .ZN(n2216) );
  INV_X1 U2032 ( .A(\REGS[4][0] ), .ZN(n538) );
  INV_X1 U2033 ( .A(\REGS[8][0] ), .ZN(n1896) );
  INV_X1 U2034 ( .A(\REGS[12][0] ), .ZN(n1960) );
  INV_X1 U2035 ( .A(\REGS[16][1] ), .ZN(n2023) );
  INV_X1 U2036 ( .A(\REGS[20][1] ), .ZN(n2087) );
  INV_X1 U2037 ( .A(\REGS[24][1] ), .ZN(n2151) );
  INV_X1 U2038 ( .A(\REGS[30][1] ), .ZN(n2215) );
  INV_X1 U2039 ( .A(\REGS[4][1] ), .ZN(n537) );
  INV_X1 U2040 ( .A(\REGS[8][1] ), .ZN(n1895) );
  INV_X1 U2041 ( .A(\REGS[12][1] ), .ZN(n1959) );
  INV_X1 U2042 ( .A(\REGS[16][2] ), .ZN(n2022) );
  INV_X1 U2043 ( .A(\REGS[20][2] ), .ZN(n2086) );
  INV_X1 U2044 ( .A(\REGS[24][2] ), .ZN(n2150) );
  INV_X1 U2045 ( .A(\REGS[30][2] ), .ZN(n2214) );
  INV_X1 U2046 ( .A(\REGS[4][2] ), .ZN(n536) );
  INV_X1 U2047 ( .A(\REGS[8][2] ), .ZN(n1894) );
  INV_X1 U2048 ( .A(\REGS[12][2] ), .ZN(n1958) );
  INV_X1 U2049 ( .A(\REGS[16][3] ), .ZN(n2021) );
  INV_X1 U2050 ( .A(\REGS[20][3] ), .ZN(n2085) );
  INV_X1 U2051 ( .A(\REGS[24][3] ), .ZN(n2149) );
  INV_X1 U2052 ( .A(\REGS[30][3] ), .ZN(n2213) );
  INV_X1 U2053 ( .A(\REGS[4][3] ), .ZN(n535) );
  INV_X1 U2054 ( .A(\REGS[8][3] ), .ZN(n1893) );
  INV_X1 U2055 ( .A(\REGS[12][3] ), .ZN(n1957) );
  INV_X1 U2056 ( .A(\REGS[16][4] ), .ZN(n2020) );
  INV_X1 U2057 ( .A(\REGS[20][4] ), .ZN(n2084) );
  INV_X1 U2058 ( .A(\REGS[24][4] ), .ZN(n2148) );
  INV_X1 U2059 ( .A(\REGS[30][4] ), .ZN(n2212) );
  INV_X1 U2060 ( .A(\REGS[4][4] ), .ZN(n534) );
  INV_X1 U2061 ( .A(\REGS[8][4] ), .ZN(n1892) );
  INV_X1 U2062 ( .A(\REGS[12][4] ), .ZN(n1956) );
  INV_X1 U2063 ( .A(\REGS[16][5] ), .ZN(n2019) );
  INV_X1 U2064 ( .A(\REGS[20][5] ), .ZN(n2083) );
  INV_X1 U2065 ( .A(\REGS[24][5] ), .ZN(n2147) );
  INV_X1 U2066 ( .A(\REGS[30][5] ), .ZN(n2211) );
  INV_X1 U2067 ( .A(\REGS[4][5] ), .ZN(n533) );
  INV_X1 U2068 ( .A(\REGS[8][5] ), .ZN(n1891) );
  INV_X1 U2069 ( .A(\REGS[12][5] ), .ZN(n1955) );
  INV_X1 U2070 ( .A(\REGS[16][6] ), .ZN(n2018) );
  INV_X1 U2071 ( .A(\REGS[20][6] ), .ZN(n2082) );
  INV_X1 U2072 ( .A(\REGS[24][6] ), .ZN(n2146) );
  INV_X1 U2073 ( .A(\REGS[30][6] ), .ZN(n2210) );
  INV_X1 U2074 ( .A(\REGS[4][6] ), .ZN(n532) );
  INV_X1 U2075 ( .A(\REGS[8][6] ), .ZN(n1890) );
  INV_X1 U2076 ( .A(\REGS[12][6] ), .ZN(n1954) );
  INV_X1 U2077 ( .A(\REGS[16][7] ), .ZN(n2017) );
  INV_X1 U2078 ( .A(\REGS[20][7] ), .ZN(n2081) );
  INV_X1 U2079 ( .A(\REGS[24][7] ), .ZN(n2145) );
  INV_X1 U2080 ( .A(\REGS[30][7] ), .ZN(n2209) );
  INV_X1 U2081 ( .A(\REGS[4][7] ), .ZN(n531) );
  INV_X1 U2082 ( .A(\REGS[8][7] ), .ZN(n1889) );
  INV_X1 U2083 ( .A(\REGS[12][7] ), .ZN(n1953) );
  INV_X1 U2084 ( .A(\REGS[16][8] ), .ZN(n2016) );
  INV_X1 U2085 ( .A(\REGS[20][8] ), .ZN(n2080) );
  INV_X1 U2086 ( .A(\REGS[24][8] ), .ZN(n2144) );
  INV_X1 U2087 ( .A(\REGS[30][8] ), .ZN(n2208) );
  INV_X1 U2088 ( .A(\REGS[4][8] ), .ZN(n530) );
  INV_X1 U2089 ( .A(\REGS[8][8] ), .ZN(n1888) );
  INV_X1 U2090 ( .A(\REGS[12][8] ), .ZN(n1952) );
  INV_X1 U2091 ( .A(\REGS[16][9] ), .ZN(n2015) );
  INV_X1 U2092 ( .A(\REGS[20][9] ), .ZN(n2079) );
  INV_X1 U2093 ( .A(\REGS[24][9] ), .ZN(n2143) );
  INV_X1 U2094 ( .A(\REGS[30][9] ), .ZN(n2207) );
  INV_X1 U2095 ( .A(\REGS[4][9] ), .ZN(n529) );
  INV_X1 U2096 ( .A(\REGS[8][9] ), .ZN(n1887) );
  INV_X1 U2097 ( .A(\REGS[12][9] ), .ZN(n1951) );
  INV_X1 U2098 ( .A(\REGS[16][10] ), .ZN(n2014) );
  INV_X1 U2099 ( .A(\REGS[20][10] ), .ZN(n2078) );
  INV_X1 U2100 ( .A(\REGS[24][10] ), .ZN(n2142) );
  INV_X1 U2101 ( .A(\REGS[30][10] ), .ZN(n2206) );
  INV_X1 U2102 ( .A(\REGS[4][10] ), .ZN(n528) );
  INV_X1 U2103 ( .A(\REGS[8][10] ), .ZN(n1886) );
  INV_X1 U2104 ( .A(\REGS[12][10] ), .ZN(n1950) );
  INV_X1 U2105 ( .A(\REGS[0][0] ), .ZN(n474) );
  INV_X1 U2106 ( .A(\REGS[0][1] ), .ZN(n473) );
  INV_X1 U2107 ( .A(\REGS[0][2] ), .ZN(n472) );
  INV_X1 U2108 ( .A(\REGS[0][3] ), .ZN(n471) );
  INV_X1 U2109 ( .A(\REGS[0][4] ), .ZN(n470) );
  INV_X1 U2110 ( .A(\REGS[0][5] ), .ZN(n469) );
  INV_X1 U2111 ( .A(\REGS[0][6] ), .ZN(n468) );
  INV_X1 U2112 ( .A(\REGS[0][7] ), .ZN(n467) );
  INV_X1 U2113 ( .A(\REGS[0][8] ), .ZN(n466) );
  INV_X1 U2114 ( .A(\REGS[0][9] ), .ZN(n465) );
  INV_X1 U2115 ( .A(\REGS[0][10] ), .ZN(n464) );
  INV_X1 U2116 ( .A(\REGS[17][0] ), .ZN(n2056) );
  INV_X1 U2117 ( .A(\REGS[21][0] ), .ZN(n2120) );
  INV_X1 U2118 ( .A(\REGS[25][0] ), .ZN(n2184) );
  INV_X1 U2119 ( .A(\REGS[31][0] ), .ZN(n2248) );
  INV_X1 U2120 ( .A(\REGS[1][0] ), .ZN(n506) );
  INV_X1 U2121 ( .A(\REGS[5][0] ), .ZN(n1864) );
  INV_X1 U2122 ( .A(\REGS[9][0] ), .ZN(n1928) );
  INV_X1 U2123 ( .A(\REGS[13][0] ), .ZN(n1992) );
  INV_X1 U2124 ( .A(\REGS[17][1] ), .ZN(n2055) );
  INV_X1 U2125 ( .A(\REGS[21][1] ), .ZN(n2119) );
  INV_X1 U2126 ( .A(\REGS[25][1] ), .ZN(n2183) );
  INV_X1 U2127 ( .A(\REGS[31][1] ), .ZN(n2247) );
  INV_X1 U2128 ( .A(\REGS[1][1] ), .ZN(n505) );
  INV_X1 U2129 ( .A(\REGS[5][1] ), .ZN(n1863) );
  INV_X1 U2130 ( .A(\REGS[9][1] ), .ZN(n1927) );
  INV_X1 U2131 ( .A(\REGS[13][1] ), .ZN(n1991) );
  INV_X1 U2132 ( .A(\REGS[17][2] ), .ZN(n2054) );
  INV_X1 U2133 ( .A(\REGS[21][2] ), .ZN(n2118) );
  INV_X1 U2134 ( .A(\REGS[25][2] ), .ZN(n2182) );
  INV_X1 U2135 ( .A(\REGS[31][2] ), .ZN(n2246) );
  INV_X1 U2136 ( .A(\REGS[1][2] ), .ZN(n504) );
  INV_X1 U2137 ( .A(\REGS[5][2] ), .ZN(n1862) );
  INV_X1 U2138 ( .A(\REGS[9][2] ), .ZN(n1926) );
  INV_X1 U2139 ( .A(\REGS[13][2] ), .ZN(n1990) );
  INV_X1 U2140 ( .A(\REGS[17][3] ), .ZN(n2053) );
  INV_X1 U2141 ( .A(\REGS[21][3] ), .ZN(n2117) );
  INV_X1 U2142 ( .A(\REGS[25][3] ), .ZN(n2181) );
  INV_X1 U2143 ( .A(\REGS[31][3] ), .ZN(n2245) );
  INV_X1 U2144 ( .A(\REGS[1][3] ), .ZN(n503) );
  INV_X1 U2145 ( .A(\REGS[5][3] ), .ZN(n1861) );
  INV_X1 U2146 ( .A(\REGS[9][3] ), .ZN(n1925) );
  INV_X1 U2147 ( .A(\REGS[13][3] ), .ZN(n1989) );
  INV_X1 U2148 ( .A(\REGS[17][4] ), .ZN(n2052) );
  INV_X1 U2149 ( .A(\REGS[21][4] ), .ZN(n2116) );
  INV_X1 U2150 ( .A(\REGS[25][4] ), .ZN(n2180) );
  INV_X1 U2151 ( .A(\REGS[31][4] ), .ZN(n2244) );
  INV_X1 U2152 ( .A(\REGS[1][4] ), .ZN(n502) );
  INV_X1 U2153 ( .A(\REGS[5][4] ), .ZN(n1860) );
  INV_X1 U2154 ( .A(\REGS[9][4] ), .ZN(n1924) );
  INV_X1 U2155 ( .A(\REGS[13][4] ), .ZN(n1988) );
  INV_X1 U2156 ( .A(\REGS[17][5] ), .ZN(n2051) );
  INV_X1 U2157 ( .A(\REGS[21][5] ), .ZN(n2115) );
  INV_X1 U2158 ( .A(\REGS[25][5] ), .ZN(n2179) );
  INV_X1 U2159 ( .A(\REGS[31][5] ), .ZN(n2243) );
  INV_X1 U2160 ( .A(\REGS[1][5] ), .ZN(n501) );
  INV_X1 U2161 ( .A(\REGS[5][5] ), .ZN(n1859) );
  INV_X1 U2162 ( .A(\REGS[9][5] ), .ZN(n1923) );
  INV_X1 U2163 ( .A(\REGS[13][5] ), .ZN(n1987) );
  INV_X1 U2164 ( .A(\REGS[17][6] ), .ZN(n2050) );
  INV_X1 U2165 ( .A(\REGS[21][6] ), .ZN(n2114) );
  INV_X1 U2166 ( .A(\REGS[25][6] ), .ZN(n2178) );
  INV_X1 U2167 ( .A(\REGS[31][6] ), .ZN(n2242) );
  INV_X1 U2168 ( .A(\REGS[1][6] ), .ZN(n500) );
  INV_X1 U2169 ( .A(\REGS[5][6] ), .ZN(n1858) );
  INV_X1 U2170 ( .A(\REGS[9][6] ), .ZN(n1922) );
  INV_X1 U2171 ( .A(\REGS[13][6] ), .ZN(n1986) );
  INV_X1 U2172 ( .A(\REGS[17][7] ), .ZN(n2049) );
  INV_X1 U2173 ( .A(\REGS[21][7] ), .ZN(n2113) );
  INV_X1 U2174 ( .A(\REGS[25][7] ), .ZN(n2177) );
  INV_X1 U2175 ( .A(\REGS[31][7] ), .ZN(n2241) );
  INV_X1 U2176 ( .A(\REGS[1][7] ), .ZN(n499) );
  INV_X1 U2177 ( .A(\REGS[5][7] ), .ZN(n1857) );
  INV_X1 U2178 ( .A(\REGS[9][7] ), .ZN(n1921) );
  INV_X1 U2179 ( .A(\REGS[13][7] ), .ZN(n1985) );
  INV_X1 U2180 ( .A(\REGS[17][8] ), .ZN(n2048) );
  INV_X1 U2181 ( .A(\REGS[21][8] ), .ZN(n2112) );
  INV_X1 U2182 ( .A(\REGS[25][8] ), .ZN(n2176) );
  INV_X1 U2183 ( .A(\REGS[31][8] ), .ZN(n2240) );
  INV_X1 U2184 ( .A(\REGS[1][8] ), .ZN(n498) );
  INV_X1 U2185 ( .A(\REGS[5][8] ), .ZN(n1856) );
  INV_X1 U2186 ( .A(\REGS[9][8] ), .ZN(n1920) );
  INV_X1 U2187 ( .A(\REGS[13][8] ), .ZN(n1984) );
  INV_X1 U2188 ( .A(\REGS[17][9] ), .ZN(n2047) );
  INV_X1 U2189 ( .A(\REGS[21][9] ), .ZN(n2111) );
  INV_X1 U2190 ( .A(\REGS[25][9] ), .ZN(n2175) );
  INV_X1 U2191 ( .A(\REGS[31][9] ), .ZN(n2239) );
  INV_X1 U2192 ( .A(\REGS[1][9] ), .ZN(n497) );
  INV_X1 U2193 ( .A(\REGS[5][9] ), .ZN(n1855) );
  INV_X1 U2194 ( .A(\REGS[9][9] ), .ZN(n1919) );
  INV_X1 U2195 ( .A(\REGS[13][9] ), .ZN(n1983) );
  INV_X1 U2196 ( .A(\REGS[17][10] ), .ZN(n2046) );
  INV_X1 U2197 ( .A(\REGS[21][10] ), .ZN(n2110) );
  INV_X1 U2198 ( .A(\REGS[25][10] ), .ZN(n2174) );
  INV_X1 U2199 ( .A(\REGS[31][10] ), .ZN(n2238) );
  INV_X1 U2200 ( .A(\REGS[1][10] ), .ZN(n496) );
  INV_X1 U2201 ( .A(\REGS[5][10] ), .ZN(n1854) );
  INV_X1 U2202 ( .A(\REGS[9][10] ), .ZN(n1918) );
  INV_X1 U2203 ( .A(\REGS[13][10] ), .ZN(n1982) );
  INV_X1 U2204 ( .A(\REGS[16][11] ), .ZN(n2013) );
  INV_X1 U2205 ( .A(\REGS[20][11] ), .ZN(n2077) );
  INV_X1 U2206 ( .A(\REGS[24][11] ), .ZN(n2141) );
  INV_X1 U2207 ( .A(\REGS[30][11] ), .ZN(n2205) );
  INV_X1 U2208 ( .A(\REGS[4][11] ), .ZN(n527) );
  INV_X1 U2209 ( .A(\REGS[8][11] ), .ZN(n1885) );
  INV_X1 U2210 ( .A(\REGS[12][11] ), .ZN(n1949) );
  INV_X1 U2211 ( .A(\REGS[16][12] ), .ZN(n2012) );
  INV_X1 U2212 ( .A(\REGS[20][12] ), .ZN(n2076) );
  INV_X1 U2213 ( .A(\REGS[24][12] ), .ZN(n2140) );
  INV_X1 U2214 ( .A(\REGS[30][12] ), .ZN(n2204) );
  INV_X1 U2215 ( .A(\REGS[4][12] ), .ZN(n526) );
  INV_X1 U2216 ( .A(\REGS[8][12] ), .ZN(n1884) );
  INV_X1 U2217 ( .A(\REGS[12][12] ), .ZN(n1948) );
  INV_X1 U2218 ( .A(\REGS[16][13] ), .ZN(n2011) );
  INV_X1 U2219 ( .A(\REGS[20][13] ), .ZN(n2075) );
  INV_X1 U2220 ( .A(\REGS[24][13] ), .ZN(n2139) );
  INV_X1 U2221 ( .A(\REGS[30][13] ), .ZN(n2203) );
  INV_X1 U2222 ( .A(\REGS[4][13] ), .ZN(n525) );
  INV_X1 U2223 ( .A(\REGS[8][13] ), .ZN(n1883) );
  INV_X1 U2224 ( .A(\REGS[12][13] ), .ZN(n1947) );
  INV_X1 U2225 ( .A(\REGS[16][14] ), .ZN(n2010) );
  INV_X1 U2226 ( .A(\REGS[20][14] ), .ZN(n2074) );
  INV_X1 U2227 ( .A(\REGS[24][14] ), .ZN(n2138) );
  INV_X1 U2228 ( .A(\REGS[30][14] ), .ZN(n2202) );
  INV_X1 U2229 ( .A(\REGS[4][14] ), .ZN(n524) );
  INV_X1 U2230 ( .A(\REGS[8][14] ), .ZN(n1882) );
  INV_X1 U2231 ( .A(\REGS[12][14] ), .ZN(n1946) );
  INV_X1 U2232 ( .A(\REGS[16][15] ), .ZN(n2009) );
  INV_X1 U2233 ( .A(\REGS[20][15] ), .ZN(n2073) );
  INV_X1 U2234 ( .A(\REGS[24][15] ), .ZN(n2137) );
  INV_X1 U2235 ( .A(\REGS[30][15] ), .ZN(n2201) );
  INV_X1 U2236 ( .A(\REGS[4][15] ), .ZN(n523) );
  INV_X1 U2237 ( .A(\REGS[8][15] ), .ZN(n1881) );
  INV_X1 U2238 ( .A(\REGS[12][15] ), .ZN(n1945) );
  INV_X1 U2239 ( .A(\REGS[16][16] ), .ZN(n2008) );
  INV_X1 U2240 ( .A(\REGS[20][16] ), .ZN(n2072) );
  INV_X1 U2241 ( .A(\REGS[24][16] ), .ZN(n2136) );
  INV_X1 U2242 ( .A(\REGS[30][16] ), .ZN(n2200) );
  INV_X1 U2243 ( .A(\REGS[4][16] ), .ZN(n522) );
  INV_X1 U2244 ( .A(\REGS[8][16] ), .ZN(n1880) );
  INV_X1 U2245 ( .A(\REGS[12][16] ), .ZN(n1944) );
  INV_X1 U2246 ( .A(\REGS[16][17] ), .ZN(n2007) );
  INV_X1 U2247 ( .A(\REGS[20][17] ), .ZN(n2071) );
  INV_X1 U2248 ( .A(\REGS[24][17] ), .ZN(n2135) );
  INV_X1 U2249 ( .A(\REGS[30][17] ), .ZN(n2199) );
  INV_X1 U2250 ( .A(\REGS[4][17] ), .ZN(n521) );
  INV_X1 U2251 ( .A(\REGS[8][17] ), .ZN(n1879) );
  INV_X1 U2252 ( .A(\REGS[12][17] ), .ZN(n1943) );
  INV_X1 U2253 ( .A(\REGS[16][18] ), .ZN(n2006) );
  INV_X1 U2254 ( .A(\REGS[20][18] ), .ZN(n2070) );
  INV_X1 U2255 ( .A(\REGS[24][18] ), .ZN(n2134) );
  INV_X1 U2256 ( .A(\REGS[30][18] ), .ZN(n2198) );
  INV_X1 U2257 ( .A(\REGS[4][18] ), .ZN(n520) );
  INV_X1 U2258 ( .A(\REGS[8][18] ), .ZN(n1878) );
  INV_X1 U2259 ( .A(\REGS[12][18] ), .ZN(n1942) );
  INV_X1 U2260 ( .A(\REGS[16][19] ), .ZN(n2005) );
  INV_X1 U2261 ( .A(\REGS[20][19] ), .ZN(n2069) );
  INV_X1 U2262 ( .A(\REGS[24][19] ), .ZN(n2133) );
  INV_X1 U2263 ( .A(\REGS[30][19] ), .ZN(n2197) );
  INV_X1 U2264 ( .A(\REGS[4][19] ), .ZN(n519) );
  INV_X1 U2265 ( .A(\REGS[8][19] ), .ZN(n1877) );
  INV_X1 U2266 ( .A(\REGS[12][19] ), .ZN(n1941) );
  INV_X1 U2267 ( .A(\REGS[16][20] ), .ZN(n2004) );
  INV_X1 U2268 ( .A(\REGS[20][20] ), .ZN(n2068) );
  INV_X1 U2269 ( .A(\REGS[24][20] ), .ZN(n2132) );
  INV_X1 U2270 ( .A(\REGS[30][20] ), .ZN(n2196) );
  INV_X1 U2271 ( .A(\REGS[4][20] ), .ZN(n518) );
  INV_X1 U2272 ( .A(\REGS[8][20] ), .ZN(n1876) );
  INV_X1 U2273 ( .A(\REGS[12][20] ), .ZN(n1940) );
  INV_X1 U2274 ( .A(\REGS[16][21] ), .ZN(n2003) );
  INV_X1 U2275 ( .A(\REGS[20][21] ), .ZN(n2067) );
  INV_X1 U2276 ( .A(\REGS[24][21] ), .ZN(n2131) );
  INV_X1 U2277 ( .A(\REGS[30][21] ), .ZN(n2195) );
  INV_X1 U2278 ( .A(\REGS[4][21] ), .ZN(n517) );
  INV_X1 U2279 ( .A(\REGS[8][21] ), .ZN(n1875) );
  INV_X1 U2280 ( .A(\REGS[12][21] ), .ZN(n1939) );
  INV_X1 U2281 ( .A(\REGS[16][22] ), .ZN(n2002) );
  INV_X1 U2282 ( .A(\REGS[20][22] ), .ZN(n2066) );
  INV_X1 U2283 ( .A(\REGS[24][22] ), .ZN(n2130) );
  INV_X1 U2284 ( .A(\REGS[30][22] ), .ZN(n2194) );
  INV_X1 U2285 ( .A(\REGS[4][22] ), .ZN(n516) );
  INV_X1 U2286 ( .A(\REGS[8][22] ), .ZN(n1874) );
  INV_X1 U2287 ( .A(\REGS[12][22] ), .ZN(n1938) );
  INV_X1 U2288 ( .A(\REGS[16][23] ), .ZN(n2001) );
  INV_X1 U2289 ( .A(\REGS[20][23] ), .ZN(n2065) );
  INV_X1 U2290 ( .A(\REGS[24][23] ), .ZN(n2129) );
  INV_X1 U2291 ( .A(\REGS[30][23] ), .ZN(n2193) );
  INV_X1 U2292 ( .A(\REGS[4][23] ), .ZN(n515) );
  INV_X1 U2293 ( .A(\REGS[8][23] ), .ZN(n1873) );
  INV_X1 U2294 ( .A(\REGS[12][23] ), .ZN(n1937) );
  INV_X1 U2295 ( .A(\REGS[16][24] ), .ZN(n2000) );
  INV_X1 U2296 ( .A(\REGS[20][24] ), .ZN(n2064) );
  INV_X1 U2297 ( .A(\REGS[24][24] ), .ZN(n2128) );
  INV_X1 U2298 ( .A(\REGS[30][24] ), .ZN(n2192) );
  INV_X1 U2299 ( .A(\REGS[4][24] ), .ZN(n514) );
  INV_X1 U2300 ( .A(\REGS[8][24] ), .ZN(n1872) );
  INV_X1 U2301 ( .A(\REGS[12][24] ), .ZN(n1936) );
  INV_X1 U2302 ( .A(\REGS[16][25] ), .ZN(n1999) );
  INV_X1 U2303 ( .A(\REGS[20][25] ), .ZN(n2063) );
  INV_X1 U2304 ( .A(\REGS[24][25] ), .ZN(n2127) );
  INV_X1 U2305 ( .A(\REGS[30][25] ), .ZN(n2191) );
  INV_X1 U2306 ( .A(\REGS[4][25] ), .ZN(n513) );
  INV_X1 U2307 ( .A(\REGS[8][25] ), .ZN(n1871) );
  INV_X1 U2308 ( .A(\REGS[12][25] ), .ZN(n1935) );
  INV_X1 U2309 ( .A(\REGS[16][26] ), .ZN(n1998) );
  INV_X1 U2310 ( .A(\REGS[20][26] ), .ZN(n2062) );
  INV_X1 U2311 ( .A(\REGS[24][26] ), .ZN(n2126) );
  INV_X1 U2312 ( .A(\REGS[30][26] ), .ZN(n2190) );
  INV_X1 U2313 ( .A(\REGS[4][26] ), .ZN(n512) );
  INV_X1 U2314 ( .A(\REGS[8][26] ), .ZN(n1870) );
  INV_X1 U2315 ( .A(\REGS[12][26] ), .ZN(n1934) );
  INV_X1 U2316 ( .A(\REGS[16][27] ), .ZN(n1997) );
  INV_X1 U2317 ( .A(\REGS[20][27] ), .ZN(n2061) );
  INV_X1 U2318 ( .A(\REGS[24][27] ), .ZN(n2125) );
  INV_X1 U2319 ( .A(\REGS[30][27] ), .ZN(n2189) );
  INV_X1 U2320 ( .A(\REGS[4][27] ), .ZN(n511) );
  INV_X1 U2321 ( .A(\REGS[8][27] ), .ZN(n1869) );
  INV_X1 U2322 ( .A(\REGS[12][27] ), .ZN(n1933) );
  INV_X1 U2323 ( .A(\REGS[16][28] ), .ZN(n1996) );
  INV_X1 U2324 ( .A(\REGS[20][28] ), .ZN(n2060) );
  INV_X1 U2325 ( .A(\REGS[24][28] ), .ZN(n2124) );
  INV_X1 U2326 ( .A(\REGS[30][28] ), .ZN(n2188) );
  INV_X1 U2327 ( .A(\REGS[4][28] ), .ZN(n510) );
  INV_X1 U2328 ( .A(\REGS[8][28] ), .ZN(n1868) );
  INV_X1 U2329 ( .A(\REGS[12][28] ), .ZN(n1932) );
  INV_X1 U2330 ( .A(\REGS[16][29] ), .ZN(n1995) );
  INV_X1 U2331 ( .A(\REGS[20][29] ), .ZN(n2059) );
  INV_X1 U2332 ( .A(\REGS[24][29] ), .ZN(n2123) );
  INV_X1 U2333 ( .A(\REGS[30][29] ), .ZN(n2187) );
  INV_X1 U2334 ( .A(\REGS[4][29] ), .ZN(n509) );
  INV_X1 U2335 ( .A(\REGS[8][29] ), .ZN(n1867) );
  INV_X1 U2336 ( .A(\REGS[12][29] ), .ZN(n1931) );
  INV_X1 U2337 ( .A(\REGS[16][30] ), .ZN(n1994) );
  INV_X1 U2338 ( .A(\REGS[20][30] ), .ZN(n2058) );
  INV_X1 U2339 ( .A(\REGS[24][30] ), .ZN(n2122) );
  INV_X1 U2340 ( .A(\REGS[30][30] ), .ZN(n2186) );
  INV_X1 U2341 ( .A(\REGS[4][30] ), .ZN(n508) );
  INV_X1 U2342 ( .A(\REGS[8][30] ), .ZN(n1866) );
  INV_X1 U2343 ( .A(\REGS[12][30] ), .ZN(n1930) );
  INV_X1 U2344 ( .A(\REGS[16][31] ), .ZN(n1993) );
  INV_X1 U2345 ( .A(\REGS[20][31] ), .ZN(n2057) );
  INV_X1 U2346 ( .A(\REGS[24][31] ), .ZN(n2121) );
  INV_X1 U2347 ( .A(\REGS[30][31] ), .ZN(n2185) );
  INV_X1 U2348 ( .A(\REGS[4][31] ), .ZN(n507) );
  INV_X1 U2349 ( .A(\REGS[8][31] ), .ZN(n1865) );
  INV_X1 U2350 ( .A(\REGS[12][31] ), .ZN(n1929) );
  INV_X1 U2351 ( .A(\REGS[0][11] ), .ZN(n463) );
  INV_X1 U2352 ( .A(\REGS[0][12] ), .ZN(n462) );
  INV_X1 U2353 ( .A(\REGS[0][13] ), .ZN(n461) );
  INV_X1 U2354 ( .A(\REGS[0][14] ), .ZN(n460) );
  INV_X1 U2355 ( .A(\REGS[0][15] ), .ZN(n459) );
  INV_X1 U2356 ( .A(\REGS[0][16] ), .ZN(n458) );
  INV_X1 U2357 ( .A(\REGS[0][17] ), .ZN(n457) );
  INV_X1 U2358 ( .A(\REGS[0][18] ), .ZN(n456) );
  INV_X1 U2359 ( .A(\REGS[0][19] ), .ZN(n455) );
  INV_X1 U2360 ( .A(\REGS[0][20] ), .ZN(n454) );
  INV_X1 U2361 ( .A(\REGS[0][21] ), .ZN(n453) );
  INV_X1 U2362 ( .A(\REGS[0][22] ), .ZN(n452) );
  INV_X1 U2363 ( .A(\REGS[0][23] ), .ZN(n451) );
  INV_X1 U2364 ( .A(\REGS[0][24] ), .ZN(n450) );
  INV_X1 U2365 ( .A(\REGS[0][25] ), .ZN(n449) );
  INV_X1 U2366 ( .A(\REGS[0][26] ), .ZN(n448) );
  INV_X1 U2367 ( .A(\REGS[0][27] ), .ZN(n447) );
  INV_X1 U2368 ( .A(\REGS[0][28] ), .ZN(n446) );
  INV_X1 U2369 ( .A(\REGS[0][29] ), .ZN(n445) );
  INV_X1 U2370 ( .A(\REGS[0][30] ), .ZN(n444) );
  INV_X1 U2371 ( .A(\REGS[0][31] ), .ZN(n443) );
  INV_X1 U2372 ( .A(ADDR_RD2[3]), .ZN(n407) );
  INV_X1 U2373 ( .A(ADDR_RD1[3]), .ZN(n403) );
  AND2_X1 U2374 ( .A1(ADDR_RD2[4]), .A2(ADDR_RD2[3]), .ZN(n1624) );
  AND2_X1 U2375 ( .A1(ADDR_RD2[4]), .A2(n407), .ZN(n1619) );
  AND2_X1 U2376 ( .A1(ADDR_RD1[4]), .A2(ADDR_RD1[3]), .ZN(n1838) );
  AND2_X1 U2377 ( .A1(ADDR_RD1[4]), .A2(n403), .ZN(n1833) );
endmodule


module MUX21_NBIT32_5 ( IN0, IN1, S, O );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] O;
  input S;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n43, n46, n47, n48, n49;

  MUX2_X2 U1 ( .A(IN1[10]), .B(IN0[10]), .S(n33), .Z(O[10]) );
  MUX2_X1 U2 ( .A(IN0[3]), .B(IN1[3]), .S(S), .Z(O[3]) );
  MUX2_X1 U3 ( .A(IN0[13]), .B(IN1[13]), .S(S), .Z(O[13]) );
  MUX2_X1 U4 ( .A(IN1[2]), .B(IN0[2]), .S(n33), .Z(O[2]) );
  MUX2_X1 U5 ( .A(IN0[4]), .B(IN1[4]), .S(S), .Z(O[4]) );
  MUX2_X1 U6 ( .A(IN0[11]), .B(IN1[11]), .S(S), .Z(O[11]) );
  MUX2_X1 U7 ( .A(IN0[14]), .B(IN1[14]), .S(S), .Z(O[14]) );
  MUX2_X1 U8 ( .A(IN0[9]), .B(IN1[9]), .S(S), .Z(O[9]) );
  MUX2_X1 U9 ( .A(IN0[7]), .B(IN1[7]), .S(S), .Z(O[7]) );
  MUX2_X1 U10 ( .A(IN0[12]), .B(IN1[12]), .S(S), .Z(O[12]) );
  MUX2_X2 U11 ( .A(IN1[1]), .B(IN0[1]), .S(n33), .Z(O[1]) );
  INV_X1 U12 ( .A(n34), .ZN(O[20]) );
  MUX2_X2 U13 ( .A(IN0[5]), .B(IN1[5]), .S(S), .Z(O[5]) );
  MUX2_X2 U14 ( .A(IN1[0]), .B(IN0[0]), .S(n33), .Z(O[0]) );
  MUX2_X2 U15 ( .A(IN0[6]), .B(IN1[6]), .S(S), .Z(O[6]) );
  MUX2_X2 U16 ( .A(IN0[8]), .B(IN1[8]), .S(S), .Z(O[8]) );
  INV_X1 U17 ( .A(n48), .ZN(O[30]) );
  AOI22_X1 U18 ( .A1(IN0[30]), .A2(n33), .B1(IN1[30]), .B2(S), .ZN(n48) );
  INV_X1 U19 ( .A(n38), .ZN(O[24]) );
  AOI22_X1 U20 ( .A1(IN0[24]), .A2(n33), .B1(IN1[24]), .B2(S), .ZN(n38) );
  INV_X1 U21 ( .A(n37), .ZN(O[23]) );
  AOI22_X1 U22 ( .A1(IN0[23]), .A2(n33), .B1(IN1[23]), .B2(S), .ZN(n37) );
  INV_X1 U23 ( .A(n39), .ZN(O[25]) );
  AOI22_X1 U24 ( .A1(IN0[25]), .A2(n33), .B1(IN1[25]), .B2(S), .ZN(n39) );
  INV_X1 U25 ( .A(n40), .ZN(O[26]) );
  AOI22_X1 U26 ( .A1(IN0[26]), .A2(n33), .B1(IN1[26]), .B2(S), .ZN(n40) );
  INV_X1 U27 ( .A(n43), .ZN(O[27]) );
  AOI22_X1 U28 ( .A1(IN0[27]), .A2(n33), .B1(IN1[27]), .B2(S), .ZN(n43) );
  AOI22_X1 U29 ( .A1(IN0[20]), .A2(n33), .B1(IN1[20]), .B2(S), .ZN(n34) );
  INV_X1 U30 ( .A(n35), .ZN(O[21]) );
  AOI22_X1 U31 ( .A1(IN0[21]), .A2(n33), .B1(IN1[21]), .B2(S), .ZN(n35) );
  INV_X1 U32 ( .A(n36), .ZN(O[22]) );
  AOI22_X1 U33 ( .A1(IN0[22]), .A2(n33), .B1(IN1[22]), .B2(S), .ZN(n36) );
  INV_X1 U34 ( .A(n49), .ZN(O[31]) );
  AOI22_X1 U35 ( .A1(IN0[31]), .A2(n33), .B1(IN1[31]), .B2(S), .ZN(n49) );
  INV_X1 U36 ( .A(n46), .ZN(O[28]) );
  AOI22_X1 U37 ( .A1(IN0[28]), .A2(n33), .B1(IN1[28]), .B2(S), .ZN(n46) );
  INV_X1 U38 ( .A(n47), .ZN(O[29]) );
  AOI22_X1 U39 ( .A1(IN0[29]), .A2(n33), .B1(IN1[29]), .B2(S), .ZN(n47) );
  MUX2_X1 U40 ( .A(IN0[15]), .B(IN1[15]), .S(S), .Z(O[15]) );
  MUX2_X1 U41 ( .A(IN0[16]), .B(IN1[16]), .S(S), .Z(O[16]) );
  MUX2_X1 U42 ( .A(IN0[17]), .B(IN1[17]), .S(S), .Z(O[17]) );
  MUX2_X1 U43 ( .A(IN0[18]), .B(IN1[18]), .S(S), .Z(O[18]) );
  MUX2_X1 U44 ( .A(IN0[19]), .B(IN1[19]), .S(S), .Z(O[19]) );
  INV_X1 U45 ( .A(S), .ZN(n33) );
endmodule


module ALU_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n233, net11615, net11613, net11612, net11524, net11523, net11522,
         net11521, net11520, net11519, net11518, net11517, net11516, net11515,
         net11514, net11513, net11511, net11505, net11502, net11501, net11500,
         net11499, net11496, net11495, net11492, net11491, net11490, net11489,
         net11486, net11485, net11482, net11481, net11480, net11479, net11476,
         net11475, net11472, net11471, net11470, net11469, net11462, net11461,
         net11460, net11459, net11456, net11455, net11450, net11449, net11448,
         net11444, net12605, net12606, net12607, net12608, net12609, net12610,
         net12611, net12614, net12615, net24602, net24601, net24626, net24672,
         net24716, net25024, net25006, net24985, net25283, n1, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232;

  AND2_X1 U1 ( .A1(n73), .A2(net11517), .ZN(net25283) );
  INV_X1 U2 ( .A(n40), .ZN(n67) );
  AND2_X1 U3 ( .A1(n45), .A2(n44), .ZN(n46) );
  NOR2_X1 U4 ( .A1(n48), .A2(n42), .ZN(n47) );
  NAND4_X1 U5 ( .A1(n43), .A2(net25006), .A3(n64), .A4(n61), .ZN(n65) );
  NOR2_X1 U6 ( .A1(n32), .A2(n33), .ZN(n52) );
  NOR2_X1 U7 ( .A1(net11520), .A2(n28), .ZN(n32) );
  NOR2_X1 U8 ( .A1(net11519), .A2(n28), .ZN(n33) );
  NOR2_X1 U9 ( .A1(n30), .A2(n27), .ZN(n51) );
  NOR2_X1 U10 ( .A1(n28), .A2(n31), .ZN(n30) );
  NOR2_X1 U11 ( .A1(n28), .A2(n29), .ZN(n27) );
  NOR2_X1 U12 ( .A1(n53), .A2(n54), .ZN(n55) );
  NAND2_X1 U13 ( .A1(net11522), .A2(net11521), .ZN(n54) );
  OAI22_X1 U14 ( .A1(net11472), .A2(n42), .B1(net11471), .B2(n42), .ZN(n53) );
  NAND2_X1 U15 ( .A1(n67), .A2(n62), .ZN(n58) );
  INV_X1 U16 ( .A(net11461), .ZN(n62) );
  NAND2_X1 U17 ( .A1(n67), .A2(n63), .ZN(n57) );
  INV_X1 U18 ( .A(net11462), .ZN(n63) );
  NOR2_X1 U19 ( .A1(n34), .A2(n36), .ZN(n59) );
  NOR2_X1 U20 ( .A1(net11524), .A2(n35), .ZN(n34) );
  NOR2_X1 U21 ( .A1(net11523), .A2(n35), .ZN(n36) );
  NAND2_X1 U22 ( .A1(n38), .A2(n39), .ZN(n35) );
  NAND2_X1 U23 ( .A1(n41), .A2(n69), .ZN(n40) );
  AND2_X1 U24 ( .A1(net11460), .A2(net11459), .ZN(n41) );
  NAND2_X1 U25 ( .A1(n4), .A2(n3), .ZN(n56) );
  AND2_X1 U26 ( .A1(n8), .A2(n156), .ZN(n134) );
  INV_X1 U27 ( .A(net24626), .ZN(n110) );
  AND2_X1 U28 ( .A1(n226), .A2(net11517), .ZN(net11490) );
  AND2_X1 U29 ( .A1(n5), .A2(n150), .ZN(n142) );
  INV_X1 U30 ( .A(net11491), .ZN(net25024) );
  AND2_X1 U31 ( .A1(net11517), .A2(net11518), .ZN(n43) );
  NAND2_X1 U32 ( .A1(net11480), .A2(net11479), .ZN(n48) );
  NOR2_X1 U33 ( .A1(net11475), .A2(n68), .ZN(n45) );
  NOR2_X1 U34 ( .A1(net11485), .A2(net11486), .ZN(n44) );
  INV_X1 U35 ( .A(net11482), .ZN(n50) );
  INV_X1 U36 ( .A(net11481), .ZN(n49) );
  NOR2_X1 U37 ( .A1(net11475), .A2(n68), .ZN(n37) );
  NAND2_X1 U38 ( .A1(net11470), .A2(net11469), .ZN(n42) );
  AND2_X1 U39 ( .A1(n154), .A2(n128), .ZN(n132) );
  NOR2_X1 U40 ( .A1(n56), .A2(n40), .ZN(n24) );
  NAND4_X1 U41 ( .A1(n57), .A2(n58), .A3(n59), .A4(n60), .ZN(n26) );
  NAND4_X1 U42 ( .A1(n51), .A2(n52), .A3(n66), .A4(n55), .ZN(n25) );
  CLKBUF_X1 U43 ( .A(n199), .Z(n1) );
  AOI21_X1 U44 ( .B1(n197), .B2(A[31]), .A(n198), .ZN(LE) );
  AOI21_X1 U45 ( .B1(n197), .B2(A[31]), .A(n198), .ZN(n233) );
  INV_X1 U46 ( .A(net24985), .ZN(n61) );
  AND2_X1 U47 ( .A1(n221), .A2(net11462), .ZN(n3) );
  OR2_X1 U48 ( .A1(n180), .A2(A[19]), .ZN(n4) );
  AND2_X1 U49 ( .A1(n3), .A2(net11522), .ZN(n5) );
  AND2_X1 U50 ( .A1(net12610), .A2(n224), .ZN(n6) );
  AND2_X1 U51 ( .A1(n71), .A2(n209), .ZN(n7) );
  AND2_X1 U52 ( .A1(net11489), .A2(n227), .ZN(n8) );
  AND2_X1 U53 ( .A1(n203), .A2(n204), .ZN(n9) );
  AND2_X1 U54 ( .A1(net11499), .A2(n231), .ZN(n10) );
  AND2_X1 U55 ( .A1(net24626), .A2(net11613), .ZN(n11) );
  AND2_X1 U56 ( .A1(net11469), .A2(n223), .ZN(n12) );
  AND2_X1 U57 ( .A1(net12605), .A2(net11514), .ZN(n13) );
  AND2_X1 U58 ( .A1(n225), .A2(net11479), .ZN(n14) );
  AND2_X1 U59 ( .A1(net11449), .A2(n219), .ZN(n15) );
  AND2_X1 U60 ( .A1(n74), .A2(net11501), .ZN(n16) );
  AND2_X1 U61 ( .A1(net25283), .A2(net11491), .ZN(n17) );
  AND2_X1 U62 ( .A1(net12615), .A2(net11524), .ZN(n18) );
  AND2_X1 U63 ( .A1(net12609), .A2(net11518), .ZN(n19) );
  AND2_X1 U64 ( .A1(net11470), .A2(net11471), .ZN(n20) );
  AOI21_X1 U65 ( .B1(n24), .B2(n25), .A(n26), .ZN(net11444) );
  INV_X1 U66 ( .A(A[3]), .ZN(n101) );
  NAND2_X1 U67 ( .A1(A[3]), .A2(n100), .ZN(net11514) );
  INV_X1 U68 ( .A(A[1]), .ZN(n99) );
  AND2_X1 U69 ( .A1(n152), .A2(n21), .ZN(n143) );
  NAND2_X1 U70 ( .A1(n215), .A2(n9), .ZN(n21) );
  NAND2_X1 U71 ( .A1(n129), .A2(n22), .ZN(n216) );
  AND2_X1 U72 ( .A1(n130), .A2(n79), .ZN(n22) );
  NAND2_X1 U73 ( .A1(n78), .A2(n79), .ZN(n23) );
  NAND2_X2 U74 ( .A1(n37), .A2(n70), .ZN(n28) );
  NAND3_X1 U75 ( .A1(net11479), .A2(n49), .A3(net11480), .ZN(n29) );
  NAND3_X1 U76 ( .A1(net11479), .A2(n50), .A3(net11480), .ZN(n31) );
  NAND3_X1 U77 ( .A1(net25024), .A2(net11489), .A3(net25283), .ZN(n64) );
  NAND3_X1 U78 ( .A1(n47), .A2(n46), .A3(n65), .ZN(n66) );
  NAND3_X1 U79 ( .A1(net11449), .A2(net11448), .A3(n71), .ZN(n60) );
  CLKBUF_X1 U80 ( .A(net11450), .Z(n71) );
  CLKBUF_X1 U81 ( .A(net11476), .Z(n68) );
  NOR2_X1 U82 ( .A1(net11455), .A2(net11456), .ZN(n39) );
  AND2_X1 U83 ( .A1(net11449), .A2(net11450), .ZN(n38) );
  AND2_X1 U84 ( .A1(n38), .A2(n39), .ZN(n69) );
  AND2_X1 U85 ( .A1(net11470), .A2(net11469), .ZN(n70) );
  AND2_X1 U86 ( .A1(net11515), .A2(net11516), .ZN(n114) );
  OR2_X1 U87 ( .A1(n193), .A2(A[6]), .ZN(n72) );
  OR2_X1 U88 ( .A1(n77), .A2(A[10]), .ZN(n73) );
  AND2_X1 U89 ( .A1(n157), .A2(n152), .ZN(n98) );
  AND2_X1 U90 ( .A1(n72), .A2(net11515), .ZN(n74) );
  AND2_X1 U91 ( .A1(n228), .A2(net11515), .ZN(net11500) );
  NAND2_X1 U92 ( .A1(net11513), .A2(net11514), .ZN(n108) );
  CLKBUF_X1 U93 ( .A(B[0]), .Z(n75) );
  AND2_X1 U94 ( .A1(n196), .A2(A[0]), .ZN(n76) );
  INV_X1 U95 ( .A(B[10]), .ZN(n77) );
  AND2_X1 U96 ( .A1(net11489), .A2(net11490), .ZN(n116) );
  AND2_X1 U97 ( .A1(net11499), .A2(net11500), .ZN(n111) );
  NOR2_X1 U98 ( .A1(net11505), .A2(n110), .ZN(n109) );
  AND2_X1 U99 ( .A1(n129), .A2(n130), .ZN(n78) );
  NOR2_X1 U100 ( .A1(n94), .A2(n144), .ZN(n79) );
  INV_X1 U101 ( .A(net11502), .ZN(n118) );
  OAI21_X1 U102 ( .B1(A[1]), .B2(n76), .A(net11613), .ZN(n104) );
  NAND2_X1 U103 ( .A1(n101), .A2(B[3]), .ZN(net24626) );
  INV_X1 U104 ( .A(B[3]), .ZN(n100) );
  INV_X1 U105 ( .A(net11501), .ZN(n117) );
  NOR2_X1 U106 ( .A1(n103), .A2(n104), .ZN(n102) );
  NAND2_X1 U107 ( .A1(n91), .A2(n82), .ZN(n80) );
  NAND2_X1 U108 ( .A1(n80), .A2(n81), .ZN(n84) );
  OR2_X1 U109 ( .A1(n164), .A2(n122), .ZN(n81) );
  AND2_X1 U110 ( .A1(n92), .A2(n83), .ZN(n82) );
  INV_X1 U111 ( .A(n164), .ZN(n83) );
  NOR2_X1 U112 ( .A1(A[1]), .A2(A[0]), .ZN(net24602) );
  OR2_X1 U113 ( .A1(n84), .A2(n85), .ZN(n86) );
  NAND2_X1 U114 ( .A1(n12), .A2(n125), .ZN(n85) );
  OAI21_X1 U115 ( .B1(net11511), .B2(n99), .A(B[1]), .ZN(n120) );
  INV_X1 U116 ( .A(n120), .ZN(n103) );
  NAND2_X1 U117 ( .A1(n86), .A2(n87), .ZN(n140) );
  OR2_X1 U118 ( .A1(n88), .A2(n127), .ZN(n87) );
  INV_X1 U119 ( .A(n125), .ZN(n88) );
  NAND2_X1 U120 ( .A1(n6), .A2(n145), .ZN(n135) );
  NAND2_X1 U121 ( .A1(n89), .A2(n90), .ZN(n91) );
  NAND2_X1 U122 ( .A1(n229), .A2(n138), .ZN(n89) );
  AND2_X1 U123 ( .A1(n137), .A2(n134), .ZN(n90) );
  NAND2_X1 U124 ( .A1(n115), .A2(n116), .ZN(n107) );
  AND3_X1 U125 ( .A1(n112), .A2(n113), .A3(n114), .ZN(n106) );
  AND2_X1 U126 ( .A1(n93), .A2(n124), .ZN(n92) );
  AND2_X2 U127 ( .A1(n224), .A2(net11519), .ZN(net11480) );
  AOI21_X1 U128 ( .B1(n105), .B2(n106), .A(n107), .ZN(net24985) );
  OAI211_X1 U129 ( .C1(n102), .C2(n108), .A(n109), .B(n111), .ZN(n105) );
  OR2_X1 U130 ( .A1(n133), .A2(n17), .ZN(n93) );
  NOR2_X1 U131 ( .A1(n162), .A2(n7), .ZN(n94) );
  NOR2_X1 U132 ( .A1(net11495), .A2(net11496), .ZN(n115) );
  INV_X1 U133 ( .A(net11492), .ZN(n119) );
  OAI211_X1 U134 ( .C1(net11615), .C2(n99), .A(net24672), .B(net24716), .ZN(
        net11612) );
  NAND2_X1 U135 ( .A1(n216), .A2(n98), .ZN(n95) );
  AND2_X1 U136 ( .A1(n95), .A2(n96), .ZN(n159) );
  OR2_X1 U137 ( .A1(n97), .A2(n9), .ZN(n96) );
  INV_X1 U138 ( .A(n152), .ZN(n97) );
  NAND3_X1 U139 ( .A1(net11499), .A2(n118), .A3(n74), .ZN(n112) );
  NAND3_X1 U140 ( .A1(net11499), .A2(n117), .A3(net11500), .ZN(n113) );
  NAND3_X1 U141 ( .A1(net11489), .A2(n119), .A3(net25283), .ZN(net25006) );
  NAND2_X1 U142 ( .A1(n140), .A2(n121), .ZN(n129) );
  AND2_X1 U143 ( .A1(n141), .A2(n132), .ZN(n121) );
  OR2_X1 U144 ( .A1(n123), .A2(n136), .ZN(n122) );
  INV_X1 U145 ( .A(n135), .ZN(n123) );
  AND2_X1 U146 ( .A1(n19), .A2(n135), .ZN(n124) );
  OR2_X1 U147 ( .A1(n126), .A2(n155), .ZN(n125) );
  INV_X1 U148 ( .A(n142), .ZN(n126) );
  AND2_X1 U149 ( .A1(n20), .A2(n142), .ZN(n127) );
  NAND2_X1 U150 ( .A1(n232), .A2(n13), .ZN(n230) );
  AND2_X1 U151 ( .A1(n15), .A2(n163), .ZN(n128) );
  OR2_X1 U152 ( .A1(n131), .A2(n18), .ZN(n130) );
  INV_X1 U153 ( .A(n128), .ZN(n131) );
  INV_X1 U154 ( .A(n156), .ZN(n133) );
  AND2_X1 U155 ( .A1(net11613), .A2(net11513), .ZN(net24716) );
  AND2_X1 U156 ( .A1(n14), .A2(n6), .ZN(n136) );
  OR2_X1 U157 ( .A1(n147), .A2(n158), .ZN(n137) );
  AND2_X1 U158 ( .A1(n16), .A2(n148), .ZN(n138) );
  AND2_X1 U159 ( .A1(n199), .A2(n146), .ZN(n139) );
  OR2_X1 U160 ( .A1(n149), .A2(n153), .ZN(n141) );
  OR2_X1 U161 ( .A1(n151), .A2(B[1]), .ZN(net24672) );
  NAND2_X1 U162 ( .A1(n168), .A2(n212), .ZN(n144) );
  NAND2_X1 U163 ( .A1(net11480), .A2(net11481), .ZN(n145) );
  OR2_X1 U164 ( .A1(B[30]), .A2(n167), .ZN(n146) );
  NAND2_X1 U165 ( .A1(n1), .A2(n146), .ZN(n197) );
  NAND2_X1 U166 ( .A1(net12607), .A2(net11516), .ZN(n147) );
  INV_X1 U167 ( .A(n147), .ZN(n148) );
  NAND2_X1 U168 ( .A1(net11460), .A2(net11461), .ZN(n149) );
  INV_X1 U169 ( .A(n149), .ZN(n150) );
  NAND2_X1 U170 ( .A1(net11612), .A2(n11), .ZN(n232) );
  INV_X1 U171 ( .A(A[0]), .ZN(net24601) );
  AND2_X1 U172 ( .A1(n75), .A2(net24601), .ZN(net11615) );
  OR2_X1 U173 ( .A1(A[30]), .A2(n160), .ZN(n152) );
  AND2_X1 U174 ( .A1(n75), .A2(net24602), .ZN(n151) );
  INV_X1 U175 ( .A(B[11]), .ZN(n188) );
  INV_X1 U176 ( .A(B[5]), .ZN(n194) );
  INV_X1 U177 ( .A(B[7]), .ZN(n192) );
  INV_X1 U178 ( .A(B[10]), .ZN(n189) );
  INV_X1 U179 ( .A(B[15]), .ZN(n184) );
  INV_X1 U180 ( .A(B[6]), .ZN(n193) );
  INV_X1 U181 ( .A(B[8]), .ZN(n191) );
  INV_X1 U182 ( .A(B[9]), .ZN(n190) );
  INV_X1 U183 ( .A(B[17]), .ZN(n182) );
  INV_X1 U184 ( .A(B[18]), .ZN(n181) );
  INV_X1 U185 ( .A(B[12]), .ZN(n187) );
  INV_X1 U186 ( .A(B[19]), .ZN(n180) );
  INV_X1 U187 ( .A(B[16]), .ZN(n183) );
  INV_X1 U188 ( .A(B[13]), .ZN(n186) );
  INV_X1 U189 ( .A(B[14]), .ZN(n185) );
  INV_X1 U190 ( .A(net11485), .ZN(net12609) );
  INV_X1 U191 ( .A(net11495), .ZN(net12607) );
  INV_X1 U192 ( .A(net11455), .ZN(net12615) );
  AND2_X1 U193 ( .A1(net11459), .A2(n221), .ZN(n153) );
  AND2_X1 U194 ( .A1(net12614), .A2(n220), .ZN(n154) );
  INV_X1 U195 ( .A(n207), .ZN(n168) );
  AND2_X1 U196 ( .A1(n4), .A2(n222), .ZN(n155) );
  AND2_X1 U197 ( .A1(net12608), .A2(n226), .ZN(n156) );
  INV_X1 U198 ( .A(B[23]), .ZN(n176) );
  INV_X1 U199 ( .A(B[27]), .ZN(n172) );
  INV_X1 U200 ( .A(net11476), .ZN(net12610) );
  INV_X1 U201 ( .A(B[24]), .ZN(n175) );
  INV_X1 U202 ( .A(B[29]), .ZN(n170) );
  INV_X1 U203 ( .A(B[25]), .ZN(n174) );
  INV_X1 U204 ( .A(B[28]), .ZN(n171) );
  INV_X1 U205 ( .A(B[26]), .ZN(n173) );
  INV_X1 U206 ( .A(B[20]), .ZN(n179) );
  INV_X1 U207 ( .A(B[21]), .ZN(n178) );
  INV_X1 U208 ( .A(B[22]), .ZN(n177) );
  INV_X1 U209 ( .A(B[0]), .ZN(n196) );
  AND2_X1 U210 ( .A1(n202), .A2(n217), .ZN(n157) );
  AND2_X1 U211 ( .A1(net12606), .A2(n72), .ZN(n158) );
  INV_X1 U212 ( .A(B[30]), .ZN(n160) );
  INV_X1 U213 ( .A(A[31]), .ZN(n166) );
  INV_X1 U214 ( .A(A[30]), .ZN(n167) );
  INV_X1 U215 ( .A(B[2]), .ZN(n161) );
  NAND2_X1 U216 ( .A1(n23), .A2(n157), .ZN(n215) );
  INV_X1 U217 ( .A(net11456), .ZN(net12614) );
  INV_X1 U218 ( .A(net11486), .ZN(net12608) );
  NAND2_X1 U219 ( .A1(n169), .A2(n218), .ZN(n162) );
  INV_X1 U220 ( .A(n162), .ZN(n163) );
  INV_X1 U221 ( .A(n208), .ZN(n169) );
  NAND2_X1 U222 ( .A1(n230), .A2(n10), .ZN(n229) );
  INV_X1 U223 ( .A(net11496), .ZN(net12606) );
  INV_X1 U224 ( .A(n213), .ZN(GE) );
  INV_X1 U225 ( .A(net11505), .ZN(net12605) );
  NAND2_X1 U226 ( .A1(net12611), .A2(net11520), .ZN(n164) );
  INV_X1 U227 ( .A(net11475), .ZN(net12611) );
  INV_X1 U228 ( .A(B[4]), .ZN(n195) );
  NAND2_X1 U229 ( .A1(n233), .A2(GE), .ZN(NE) );
  AOI21_X1 U230 ( .B1(n139), .B2(n166), .A(B[31]), .ZN(n198) );
  OAI211_X1 U231 ( .C1(n200), .C2(n201), .A(n202), .B(n203), .ZN(n199) );
  NAND2_X1 U232 ( .A1(n204), .A2(n205), .ZN(n201) );
  AOI211_X1 U233 ( .C1(net11444), .C2(n206), .A(n207), .B(n208), .ZN(n200) );
  NAND2_X1 U234 ( .A1(n209), .A2(n210), .ZN(net11448) );
  NAND2_X1 U235 ( .A1(n196), .A2(A[0]), .ZN(net11511) );
  AND2_X1 U236 ( .A1(n211), .A2(n212), .ZN(n206) );
  OAI21_X1 U237 ( .B1(n143), .B2(A[31]), .A(n214), .ZN(n213) );
  OAI21_X1 U238 ( .B1(n159), .B2(n166), .A(B[31]), .ZN(n214) );
  XOR2_X1 U239 ( .A(n167), .B(B[30]), .Z(n203) );
  NAND2_X1 U240 ( .A1(A[29]), .A2(n170), .ZN(n204) );
  OR2_X1 U241 ( .A1(n170), .A2(A[29]), .ZN(n202) );
  NAND2_X1 U242 ( .A1(n217), .A2(n205), .ZN(n207) );
  NAND2_X1 U243 ( .A1(A[28]), .A2(n171), .ZN(n205) );
  OR2_X1 U244 ( .A1(n171), .A2(A[28]), .ZN(n217) );
  NAND2_X1 U245 ( .A1(A[27]), .A2(n172), .ZN(n212) );
  NOR2_X1 U246 ( .A1(n172), .A2(A[27]), .ZN(n208) );
  AND2_X1 U247 ( .A1(n218), .A2(n211), .ZN(net11450) );
  NAND2_X1 U248 ( .A1(A[26]), .A2(n173), .ZN(n211) );
  OR2_X1 U249 ( .A1(n173), .A2(A[26]), .ZN(n218) );
  NAND2_X1 U250 ( .A1(A[25]), .A2(n174), .ZN(n209) );
  OR2_X1 U251 ( .A1(n174), .A2(A[25]), .ZN(net11449) );
  NAND2_X1 U252 ( .A1(n219), .A2(n210), .ZN(net11455) );
  NAND2_X1 U253 ( .A1(A[24]), .A2(n175), .ZN(n210) );
  OR2_X1 U254 ( .A1(n175), .A2(A[24]), .ZN(n219) );
  NAND2_X1 U255 ( .A1(A[23]), .A2(n176), .ZN(net11524) );
  NOR2_X1 U256 ( .A1(n176), .A2(A[23]), .ZN(net11456) );
  AND2_X1 U257 ( .A1(n220), .A2(net11523), .ZN(net11460) );
  NAND2_X1 U258 ( .A1(A[22]), .A2(n177), .ZN(net11523) );
  OR2_X1 U259 ( .A1(n177), .A2(A[22]), .ZN(n220) );
  NAND2_X1 U260 ( .A1(A[21]), .A2(n178), .ZN(net11461) );
  OR2_X1 U261 ( .A1(n178), .A2(A[21]), .ZN(net11459) );
  NAND2_X1 U262 ( .A1(A[20]), .A2(n179), .ZN(net11462) );
  OR2_X1 U263 ( .A1(n179), .A2(A[20]), .ZN(n221) );
  NAND2_X1 U264 ( .A1(A[19]), .A2(n180), .ZN(net11522) );
  AND2_X1 U265 ( .A1(n222), .A2(net11521), .ZN(net11470) );
  NAND2_X1 U266 ( .A1(A[18]), .A2(n181), .ZN(net11521) );
  OR2_X1 U267 ( .A1(n181), .A2(A[18]), .ZN(n222) );
  NAND2_X1 U268 ( .A1(A[17]), .A2(n182), .ZN(net11471) );
  OR2_X1 U269 ( .A1(n182), .A2(A[17]), .ZN(net11469) );
  NAND2_X1 U270 ( .A1(n223), .A2(net11472), .ZN(net11475) );
  NAND2_X1 U271 ( .A1(A[16]), .A2(n183), .ZN(net11472) );
  OR2_X1 U272 ( .A1(n183), .A2(A[16]), .ZN(n223) );
  NAND2_X1 U273 ( .A1(A[15]), .A2(n184), .ZN(net11520) );
  NOR2_X1 U274 ( .A1(n184), .A2(A[15]), .ZN(net11476) );
  NAND2_X1 U275 ( .A1(A[14]), .A2(n185), .ZN(net11519) );
  OR2_X1 U276 ( .A1(n185), .A2(A[14]), .ZN(n224) );
  NAND2_X1 U277 ( .A1(A[13]), .A2(n186), .ZN(net11481) );
  OR2_X1 U278 ( .A1(n186), .A2(A[13]), .ZN(net11479) );
  NAND2_X1 U279 ( .A1(n225), .A2(net11482), .ZN(net11485) );
  NAND2_X1 U280 ( .A1(A[12]), .A2(n187), .ZN(net11482) );
  OR2_X1 U281 ( .A1(n187), .A2(A[12]), .ZN(n225) );
  NAND2_X1 U282 ( .A1(A[11]), .A2(n188), .ZN(net11518) );
  NOR2_X1 U283 ( .A1(n188), .A2(A[11]), .ZN(net11486) );
  NAND2_X1 U284 ( .A1(A[10]), .A2(n189), .ZN(net11517) );
  OR2_X1 U285 ( .A1(n77), .A2(A[10]), .ZN(n226) );
  NAND2_X1 U286 ( .A1(A[9]), .A2(n190), .ZN(net11491) );
  OR2_X1 U287 ( .A1(n190), .A2(A[9]), .ZN(net11489) );
  NAND2_X1 U288 ( .A1(n227), .A2(net11492), .ZN(net11495) );
  NAND2_X1 U289 ( .A1(A[8]), .A2(n191), .ZN(net11492) );
  OR2_X1 U290 ( .A1(n191), .A2(A[8]), .ZN(n227) );
  NAND2_X1 U291 ( .A1(A[7]), .A2(n192), .ZN(net11516) );
  NOR2_X1 U292 ( .A1(n192), .A2(A[7]), .ZN(net11496) );
  NAND2_X1 U293 ( .A1(A[6]), .A2(n193), .ZN(net11515) );
  OR2_X1 U294 ( .A1(n193), .A2(A[6]), .ZN(n228) );
  NAND2_X1 U295 ( .A1(A[5]), .A2(n194), .ZN(net11501) );
  OR2_X1 U296 ( .A1(n194), .A2(A[5]), .ZN(net11499) );
  NAND2_X1 U297 ( .A1(n231), .A2(net11502), .ZN(net11505) );
  NAND2_X1 U298 ( .A1(A[4]), .A2(n195), .ZN(net11502) );
  OR2_X1 U299 ( .A1(n195), .A2(A[4]), .ZN(n231) );
  NAND2_X1 U300 ( .A1(n161), .A2(A[2]), .ZN(net11513) );
  OR2_X1 U301 ( .A1(n161), .A2(A[2]), .ZN(net11613) );
endmodule


module ALU_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   net15501, net15500, net15499, net15496, net15491, net15475, net15471,
         net15463, net15462, net15460, net15458, net15451, net15429, net15428,
         net24577, net25175, net25215, net25247, net25312, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285;

  INV_X1 U3 ( .A(B[27]), .ZN(n98) );
  NAND2_X1 U4 ( .A1(n15), .A2(B[29]), .ZN(n5) );
  INV_X1 U5 ( .A(A[29]), .ZN(n15) );
  INV_X1 U6 ( .A(B[29]), .ZN(n16) );
  NOR2_X1 U7 ( .A1(net15462), .A2(n9), .ZN(n13) );
  INV_X1 U8 ( .A(net15463), .ZN(n11) );
  NAND2_X1 U9 ( .A1(A[28]), .A2(n19), .ZN(n20) );
  INV_X1 U10 ( .A(B[28]), .ZN(n19) );
  INV_X1 U11 ( .A(A[30]), .ZN(n10) );
  INV_X1 U12 ( .A(net15491), .ZN(n9) );
  AND4_X1 U13 ( .A1(n71), .A2(n64), .A3(n58), .A4(n56), .ZN(n33) );
  NOR2_X1 U14 ( .A1(B[30]), .A2(n10), .ZN(n17) );
  NAND2_X1 U15 ( .A1(B[30]), .A2(n10), .ZN(n22) );
  NAND2_X1 U16 ( .A1(A[29]), .A2(n16), .ZN(n8) );
  NAND2_X1 U17 ( .A1(n5), .A2(n6), .ZN(net24577) );
  NAND2_X1 U18 ( .A1(A[29]), .A2(n16), .ZN(n6) );
  INV_X1 U19 ( .A(n20), .ZN(net15458) );
  NAND2_X1 U20 ( .A1(net15475), .A2(net15491), .ZN(net15496) );
  AND2_X1 U21 ( .A1(B[28]), .A2(net15460), .ZN(n1) );
  AND4_X1 U22 ( .A1(n235), .A2(n239), .A3(n48), .A4(n53), .ZN(n2) );
  XOR2_X1 U23 ( .A(A[30]), .B(B[30]), .Z(n3) );
  NAND2_X1 U24 ( .A1(A[2]), .A2(n280), .ZN(n4) );
  OAI21_X1 U25 ( .B1(n12), .B2(n1), .A(n20), .ZN(n21) );
  NAND2_X1 U26 ( .A1(n21), .A2(n5), .ZN(n7) );
  INV_X1 U27 ( .A(n21), .ZN(net25175) );
  AOI21_X1 U28 ( .B1(n13), .B2(n14), .A(n11), .ZN(n12) );
  OAI21_X1 U29 ( .B1(net15500), .B2(net15499), .A(net15501), .ZN(n14) );
  OAI21_X1 U30 ( .B1(net15429), .B2(n17), .A(n22), .ZN(n18) );
  XNOR2_X1 U31 ( .A(net15428), .B(n18), .ZN(DIFF[31]) );
  NAND2_X1 U32 ( .A1(net25312), .A2(net15491), .ZN(net25247) );
  NAND2_X1 U33 ( .A1(n7), .A2(n8), .ZN(net15429) );
  OAI21_X1 U34 ( .B1(net25247), .B2(net15462), .A(net15463), .ZN(net15451) );
  BUF_X1 U35 ( .A(n84), .Z(n23) );
  AND2_X1 U36 ( .A1(A[2]), .A2(n280), .ZN(n30) );
  NAND4_X1 U37 ( .A1(n235), .A2(n239), .A3(n48), .A4(n53), .ZN(n24) );
  AND2_X1 U38 ( .A1(n271), .A2(n272), .ZN(n25) );
  CLKBUF_X1 U39 ( .A(n35), .Z(n26) );
  AND2_X1 U40 ( .A1(n264), .A2(A[6]), .ZN(n35) );
  CLKBUF_X1 U41 ( .A(n206), .Z(n27) );
  CLKBUF_X1 U42 ( .A(n58), .Z(n28) );
  CLKBUF_X1 U43 ( .A(n36), .Z(n29) );
  OAI21_X1 U44 ( .B1(net15499), .B2(net15500), .A(net15501), .ZN(net25312) );
  CLKBUF_X1 U45 ( .A(n161), .Z(n31) );
  OAI21_X2 U46 ( .B1(n69), .B2(n203), .A(n256), .ZN(n51) );
  CLKBUF_X1 U47 ( .A(n142), .Z(n32) );
  CLKBUF_X1 U48 ( .A(n106), .Z(n34) );
  CLKBUF_X1 U49 ( .A(net15499), .Z(net25215) );
  INV_X1 U50 ( .A(n29), .ZN(n162) );
  XNOR2_X1 U51 ( .A(net15429), .B(n3), .ZN(DIFF[30]) );
  INV_X1 U52 ( .A(n26), .ZN(n66) );
  AND2_X1 U53 ( .A1(B[0]), .A2(n284), .ZN(n36) );
  CLKBUF_X1 U54 ( .A(n70), .Z(n37) );
  OAI21_X1 U55 ( .B1(n32), .B2(n143), .A(n144), .ZN(n38) );
  NAND2_X1 U56 ( .A1(A[1]), .A2(n276), .ZN(n39) );
  NAND2_X1 U57 ( .A1(A[1]), .A2(n276), .ZN(n40) );
  CLKBUF_X1 U58 ( .A(n175), .Z(n41) );
  XOR2_X1 U59 ( .A(n42), .B(n226), .Z(DIFF[12]) );
  AND2_X1 U60 ( .A1(n199), .A2(n207), .ZN(n42) );
  XOR2_X1 U61 ( .A(net15451), .B(n43), .Z(DIFF[28]) );
  NOR2_X1 U62 ( .A1(n1), .A2(net15458), .ZN(n43) );
  XOR2_X1 U63 ( .A(net25175), .B(net24577), .Z(DIFF[29]) );
  XOR2_X1 U64 ( .A(n54), .B(n55), .Z(DIFF[7]) );
  OAI21_X1 U65 ( .B1(n229), .B2(n24), .A(n230), .ZN(n226) );
  NOR2_X1 U66 ( .A1(n24), .A2(n202), .ZN(n205) );
  NOR2_X1 U67 ( .A1(n202), .A2(n187), .ZN(n201) );
  NAND2_X1 U68 ( .A1(n25), .A2(n186), .ZN(n73) );
  NAND4_X1 U69 ( .A1(n235), .A2(n239), .A3(n48), .A4(n53), .ZN(n187) );
  OAI21_X1 U70 ( .B1(n61), .B2(n62), .A(n63), .ZN(n59) );
  OAI21_X1 U71 ( .B1(n218), .B2(n219), .A(n198), .ZN(n214) );
  NAND4_X1 U72 ( .A1(n207), .A2(n196), .A3(n208), .A4(n188), .ZN(n202) );
  OAI21_X1 U73 ( .B1(n142), .B2(n143), .A(n144), .ZN(n137) );
  AOI21_X1 U74 ( .B1(n145), .B2(n146), .A(n147), .ZN(n144) );
  OAI21_X1 U75 ( .B1(n231), .B2(n232), .A(n233), .ZN(n204) );
  NAND2_X1 U76 ( .A1(n235), .A2(n48), .ZN(n232) );
  AOI21_X1 U77 ( .B1(n234), .B2(n235), .A(n236), .ZN(n233) );
  NAND2_X1 U78 ( .A1(n239), .A2(n240), .ZN(n231) );
  AOI21_X1 U79 ( .B1(n86), .B2(n87), .A(n45), .ZN(net15463) );
  OAI21_X1 U80 ( .B1(n88), .B2(n89), .A(n90), .ZN(n87) );
  OAI21_X1 U81 ( .B1(net25215), .B2(net15500), .A(net15501), .ZN(n108) );
  AOI21_X1 U82 ( .B1(n113), .B2(n114), .A(n115), .ZN(net15501) );
  NAND4_X1 U83 ( .A1(n180), .A2(n183), .A3(n181), .A4(n182), .ZN(n175) );
  AOI21_X1 U84 ( .B1(n188), .B2(n189), .A(n190), .ZN(n182) );
  AOI22_X1 U85 ( .A1(n184), .A2(n204), .B1(n206), .B2(n205), .ZN(n180) );
  OAI21_X1 U86 ( .B1(n224), .B2(n225), .A(n199), .ZN(n220) );
  OAI21_X1 U87 ( .B1(n68), .B2(n69), .A(n37), .ZN(n65) );
  OAI21_X1 U88 ( .B1(n251), .B2(n46), .A(n49), .ZN(n247) );
  NAND4_X1 U89 ( .A1(n71), .A2(n64), .A3(n28), .A4(n56), .ZN(n203) );
  NAND2_X1 U90 ( .A1(n156), .A2(n176), .ZN(n179) );
  NAND2_X1 U91 ( .A1(n148), .A2(n145), .ZN(n163) );
  NAND2_X1 U92 ( .A1(n124), .A2(n138), .ZN(n141) );
  NAND2_X1 U93 ( .A1(n198), .A2(n196), .ZN(n223) );
  XOR2_X1 U94 ( .A(n128), .B(n131), .Z(DIFF[22]) );
  NAND2_X1 U95 ( .A1(n119), .A2(n125), .ZN(n131) );
  NAND2_X1 U96 ( .A1(n52), .A2(n53), .ZN(n50) );
  XOR2_X1 U97 ( .A(n44), .B(n74), .Z(DIFF[3]) );
  AND2_X1 U98 ( .A1(n79), .A2(n80), .ZN(n44) );
  NAND2_X1 U99 ( .A1(n64), .A2(n63), .ZN(n67) );
  NAND2_X1 U100 ( .A1(n238), .A2(n239), .ZN(n250) );
  NAND2_X1 U101 ( .A1(n237), .A2(n235), .ZN(n243) );
  OAI21_X1 U102 ( .B1(n245), .B2(n246), .A(n238), .ZN(n244) );
  XOR2_X1 U103 ( .A(n46), .B(n47), .Z(DIFF[9]) );
  NAND2_X1 U104 ( .A1(n48), .A2(n49), .ZN(n47) );
  OAI21_X1 U105 ( .B1(n192), .B2(n193), .A(n194), .ZN(n189) );
  AOI21_X1 U106 ( .B1(n195), .B2(n196), .A(n197), .ZN(n192) );
  OAI21_X1 U107 ( .B1(n117), .B2(n118), .A(n119), .ZN(n114) );
  AOI21_X1 U108 ( .B1(n120), .B2(n121), .A(n122), .ZN(n117) );
  NAND2_X1 U109 ( .A1(net25215), .A2(n124), .ZN(n135) );
  NAND2_X1 U110 ( .A1(n32), .A2(n156), .ZN(n171) );
  NAND2_X1 U111 ( .A1(n257), .A2(n258), .ZN(n206) );
  AOI21_X1 U112 ( .B1(n35), .B2(n56), .A(n262), .ZN(n257) );
  NAND4_X1 U113 ( .A1(n259), .A2(n64), .A3(n58), .A4(n56), .ZN(n258) );
  NAND2_X1 U114 ( .A1(n29), .A2(n31), .ZN(n85) );
  NAND2_X1 U115 ( .A1(n105), .A2(n94), .ZN(n100) );
  NAND2_X1 U116 ( .A1(n92), .A2(n106), .ZN(n105) );
  OAI21_X1 U117 ( .B1(n128), .B2(n118), .A(n119), .ZN(n127) );
  NAND2_X1 U118 ( .A1(net25247), .A2(net15475), .ZN(n106) );
  NAND2_X1 U119 ( .A1(n170), .A2(n155), .ZN(n166) );
  NAND2_X1 U120 ( .A1(n153), .A2(n171), .ZN(n170) );
  NAND2_X1 U121 ( .A1(n82), .A2(n39), .ZN(n78) );
  NAND2_X1 U122 ( .A1(n23), .A2(n85), .ZN(n82) );
  XNOR2_X1 U123 ( .A(n81), .B(n78), .ZN(DIFF[2]) );
  NAND2_X1 U124 ( .A1(n77), .A2(n4), .ZN(n81) );
  XNOR2_X1 U125 ( .A(n100), .B(n102), .ZN(DIFF[26]) );
  NAND2_X1 U126 ( .A1(n90), .A2(n91), .ZN(n102) );
  AOI21_X1 U127 ( .B1(n28), .B2(n59), .A(n26), .ZN(n54) );
  NAND2_X1 U128 ( .A1(n56), .A2(n57), .ZN(n55) );
  XNOR2_X1 U129 ( .A(n60), .B(n59), .ZN(DIFF[6]) );
  NAND2_X1 U130 ( .A1(n28), .A2(n66), .ZN(n60) );
  XNOR2_X1 U131 ( .A(n217), .B(n214), .ZN(DIFF[14]) );
  NAND2_X1 U132 ( .A1(n194), .A2(n208), .ZN(n217) );
  XNOR2_X1 U133 ( .A(n174), .B(n171), .ZN(DIFF[17]) );
  NAND2_X1 U134 ( .A1(n155), .A2(n153), .ZN(n174) );
  XNOR2_X1 U135 ( .A(n107), .B(n34), .ZN(DIFF[25]) );
  NAND2_X1 U136 ( .A1(n94), .A2(n92), .ZN(n107) );
  XNOR2_X1 U137 ( .A(n95), .B(n96), .ZN(DIFF[27]) );
  AOI21_X1 U138 ( .B1(n91), .B2(n100), .A(n101), .ZN(n95) );
  XNOR2_X1 U139 ( .A(n169), .B(n166), .ZN(DIFF[18]) );
  NAND2_X1 U140 ( .A1(n151), .A2(n157), .ZN(n169) );
  XNOR2_X1 U141 ( .A(n136), .B(n135), .ZN(DIFF[21]) );
  NAND2_X1 U142 ( .A1(n123), .A2(n121), .ZN(n136) );
  XNOR2_X1 U143 ( .A(n72), .B(n73), .ZN(DIFF[4]) );
  NAND2_X1 U144 ( .A1(n37), .A2(n71), .ZN(n72) );
  XNOR2_X1 U145 ( .A(n108), .B(net15496), .ZN(DIFF[24]) );
  XNOR2_X1 U146 ( .A(n160), .B(n85), .ZN(DIFF[1]) );
  NAND2_X1 U147 ( .A1(n23), .A2(n40), .ZN(n160) );
  NAND2_X1 U148 ( .A1(n175), .A2(n176), .ZN(n142) );
  AOI21_X1 U149 ( .B1(net15471), .B2(n92), .A(n93), .ZN(n88) );
  OAI21_X1 U150 ( .B1(n149), .B2(n150), .A(n151), .ZN(n146) );
  AOI21_X1 U151 ( .B1(n152), .B2(n153), .A(n154), .ZN(n149) );
  NAND2_X1 U152 ( .A1(n137), .A2(n138), .ZN(net15499) );
  NAND2_X1 U153 ( .A1(n49), .A2(n52), .ZN(n240) );
  NAND2_X1 U154 ( .A1(n70), .A2(n63), .ZN(n259) );
  NAND2_X1 U155 ( .A1(n83), .A2(n161), .ZN(n273) );
  AND2_X1 U156 ( .A1(n134), .A2(n123), .ZN(n128) );
  NAND2_X1 U157 ( .A1(n121), .A2(n135), .ZN(n134) );
  NAND2_X1 U158 ( .A1(n271), .A2(n272), .ZN(n200) );
  AOI21_X1 U159 ( .B1(n30), .B2(n79), .A(n277), .ZN(n271) );
  NAND4_X1 U160 ( .A1(n273), .A2(n23), .A3(n77), .A4(n79), .ZN(n272) );
  AND2_X1 U161 ( .A1(n253), .A2(n52), .ZN(n46) );
  NAND2_X1 U162 ( .A1(n51), .A2(n53), .ZN(n253) );
  XNOR2_X1 U163 ( .A(n211), .B(n212), .ZN(DIFF[15]) );
  NAND2_X1 U164 ( .A1(n191), .A2(n188), .ZN(n211) );
  OAI21_X1 U165 ( .B1(n213), .B2(n193), .A(n194), .ZN(n212) );
  NAND2_X1 U166 ( .A1(n31), .A2(n162), .ZN(DIFF[0]) );
  NAND2_X1 U167 ( .A1(n116), .A2(n113), .ZN(n126) );
  INV_X1 U168 ( .A(A[2]), .ZN(n274) );
  NAND2_X1 U169 ( .A1(A[9]), .A2(n252), .ZN(n49) );
  INV_X1 U170 ( .A(B[9]), .ZN(n252) );
  NAND2_X1 U171 ( .A1(B[11]), .A2(n248), .ZN(n235) );
  INV_X1 U172 ( .A(A[11]), .ZN(n248) );
  NAND2_X1 U173 ( .A1(B[7]), .A2(n265), .ZN(n56) );
  INV_X1 U174 ( .A(A[7]), .ZN(n265) );
  NAND2_X1 U175 ( .A1(A[26]), .A2(n104), .ZN(n90) );
  INV_X1 U176 ( .A(B[26]), .ZN(n104) );
  NAND2_X1 U177 ( .A1(A[22]), .A2(n133), .ZN(n119) );
  INV_X1 U178 ( .A(B[22]), .ZN(n133) );
  NAND2_X1 U179 ( .A1(A[14]), .A2(n222), .ZN(n194) );
  INV_X1 U180 ( .A(B[14]), .ZN(n222) );
  NAND2_X1 U181 ( .A1(A[5]), .A2(n261), .ZN(n63) );
  INV_X1 U182 ( .A(B[5]), .ZN(n261) );
  NAND2_X1 U183 ( .A1(B[6]), .A2(n266), .ZN(n58) );
  INV_X1 U184 ( .A(A[6]), .ZN(n266) );
  INV_X1 U185 ( .A(A[4]), .ZN(n268) );
  NAND2_X1 U186 ( .A1(A[4]), .A2(n260), .ZN(n70) );
  NAND2_X1 U187 ( .A1(A[25]), .A2(n110), .ZN(n94) );
  INV_X1 U188 ( .A(B[25]), .ZN(n110) );
  NAND2_X1 U189 ( .A1(A[16]), .A2(n210), .ZN(n156) );
  INV_X1 U190 ( .A(B[16]), .ZN(n210) );
  INV_X1 U191 ( .A(A[0]), .ZN(n284) );
  NAND2_X1 U192 ( .A1(A[12]), .A2(n242), .ZN(n199) );
  INV_X1 U193 ( .A(B[12]), .ZN(n242) );
  NAND2_X1 U194 ( .A1(A[13]), .A2(n228), .ZN(n198) );
  INV_X1 U195 ( .A(B[13]), .ZN(n228) );
  NAND2_X1 U196 ( .A1(B[9]), .A2(n281), .ZN(n48) );
  INV_X1 U197 ( .A(A[9]), .ZN(n281) );
  NAND2_X1 U198 ( .A1(A[7]), .A2(n263), .ZN(n57) );
  INV_X1 U199 ( .A(B[7]), .ZN(n263) );
  NAND2_X1 U200 ( .A1(A[3]), .A2(n278), .ZN(n80) );
  NAND2_X1 U201 ( .A1(B[17]), .A2(n177), .ZN(n153) );
  INV_X1 U202 ( .A(A[17]), .ZN(n177) );
  NAND2_X1 U203 ( .A1(B[15]), .A2(n215), .ZN(n188) );
  INV_X1 U204 ( .A(A[15]), .ZN(n215) );
  NAND2_X1 U205 ( .A1(A[15]), .A2(n216), .ZN(n191) );
  INV_X1 U206 ( .A(B[15]), .ZN(n216) );
  NAND2_X1 U207 ( .A1(B[14]), .A2(n221), .ZN(n208) );
  INV_X1 U208 ( .A(A[14]), .ZN(n221) );
  NAND2_X1 U209 ( .A1(B[12]), .A2(n241), .ZN(n207) );
  INV_X1 U210 ( .A(A[12]), .ZN(n241) );
  NAND2_X1 U211 ( .A1(A[24]), .A2(n112), .ZN(net15475) );
  INV_X1 U212 ( .A(B[24]), .ZN(n112) );
  NAND2_X1 U213 ( .A1(B[18]), .A2(n172), .ZN(n157) );
  INV_X1 U214 ( .A(A[18]), .ZN(n172) );
  NAND2_X1 U215 ( .A1(B[16]), .A2(n209), .ZN(n176) );
  INV_X1 U216 ( .A(A[16]), .ZN(n209) );
  NAND2_X1 U217 ( .A1(A[23]), .A2(n130), .ZN(n116) );
  INV_X1 U218 ( .A(B[23]), .ZN(n130) );
  NAND2_X1 U219 ( .A1(B[21]), .A2(n139), .ZN(n121) );
  INV_X1 U220 ( .A(A[21]), .ZN(n139) );
  NAND2_X1 U221 ( .A1(B[25]), .A2(n109), .ZN(n92) );
  INV_X1 U222 ( .A(A[25]), .ZN(n109) );
  NAND2_X1 U223 ( .A1(B[1]), .A2(n275), .ZN(n84) );
  INV_X1 U224 ( .A(A[1]), .ZN(n275) );
  NAND2_X1 U225 ( .A1(B[19]), .A2(n167), .ZN(n145) );
  INV_X1 U226 ( .A(A[19]), .ZN(n167) );
  NAND2_X1 U227 ( .A1(B[26]), .A2(n103), .ZN(n91) );
  INV_X1 U228 ( .A(A[26]), .ZN(n103) );
  NAND2_X1 U229 ( .A1(B[10]), .A2(n282), .ZN(n239) );
  INV_X1 U230 ( .A(A[10]), .ZN(n282) );
  NAND2_X1 U231 ( .A1(B[8]), .A2(n255), .ZN(n53) );
  INV_X1 U232 ( .A(A[8]), .ZN(n255) );
  NAND2_X1 U233 ( .A1(A[0]), .A2(n285), .ZN(n161) );
  INV_X1 U234 ( .A(B[0]), .ZN(n285) );
  INV_X1 U235 ( .A(A[3]), .ZN(n279) );
  NAND2_X1 U236 ( .A1(B[13]), .A2(n227), .ZN(n196) );
  INV_X1 U237 ( .A(A[13]), .ZN(n227) );
  NAND2_X1 U238 ( .A1(B[5]), .A2(n267), .ZN(n64) );
  INV_X1 U239 ( .A(A[5]), .ZN(n267) );
  NAND2_X1 U240 ( .A1(B[23]), .A2(n129), .ZN(n113) );
  INV_X1 U241 ( .A(A[23]), .ZN(n129) );
  AND2_X1 U242 ( .A1(A[27]), .A2(n98), .ZN(n45) );
  NAND2_X1 U243 ( .A1(A[11]), .A2(n249), .ZN(n237) );
  INV_X1 U244 ( .A(B[11]), .ZN(n249) );
  XNOR2_X1 U245 ( .A(B[31]), .B(A[31]), .ZN(net15428) );
  NAND2_X1 U246 ( .A1(A[10]), .A2(n283), .ZN(n238) );
  INV_X1 U247 ( .A(B[10]), .ZN(n283) );
  NAND2_X1 U248 ( .A1(B[24]), .A2(n111), .ZN(net15491) );
  INV_X1 U249 ( .A(A[24]), .ZN(n111) );
  NAND2_X1 U250 ( .A1(B[20]), .A2(n158), .ZN(n138) );
  INV_X1 U251 ( .A(A[20]), .ZN(n158) );
  NAND2_X1 U252 ( .A1(B[27]), .A2(n99), .ZN(n86) );
  INV_X1 U253 ( .A(A[27]), .ZN(n99) );
  INV_X1 U254 ( .A(B[6]), .ZN(n264) );
  NAND2_X1 U255 ( .A1(A[8]), .A2(n254), .ZN(n52) );
  INV_X1 U256 ( .A(B[8]), .ZN(n254) );
  NAND2_X1 U257 ( .A1(B[22]), .A2(n132), .ZN(n125) );
  INV_X1 U258 ( .A(A[22]), .ZN(n132) );
  NAND2_X1 U259 ( .A1(A[17]), .A2(n178), .ZN(n155) );
  INV_X1 U260 ( .A(B[17]), .ZN(n178) );
  NAND2_X1 U261 ( .A1(A[18]), .A2(n173), .ZN(n151) );
  INV_X1 U262 ( .A(B[18]), .ZN(n173) );
  INV_X1 U263 ( .A(A[28]), .ZN(net15460) );
  NAND2_X1 U264 ( .A1(A[19]), .A2(n168), .ZN(n148) );
  INV_X1 U265 ( .A(B[19]), .ZN(n168) );
  NAND2_X1 U266 ( .A1(A[1]), .A2(n276), .ZN(n83) );
  INV_X1 U267 ( .A(B[1]), .ZN(n276) );
  NAND2_X1 U268 ( .A1(A[20]), .A2(n159), .ZN(n124) );
  INV_X1 U269 ( .A(B[20]), .ZN(n159) );
  NAND2_X1 U270 ( .A1(A[21]), .A2(n140), .ZN(n123) );
  INV_X1 U271 ( .A(B[21]), .ZN(n140) );
  NAND2_X1 U272 ( .A1(B[3]), .A2(n279), .ZN(n79) );
  INV_X1 U273 ( .A(B[3]), .ZN(n278) );
  NAND2_X1 U274 ( .A1(B[4]), .A2(n268), .ZN(n71) );
  INV_X1 U275 ( .A(B[4]), .ZN(n260) );
  INV_X1 U276 ( .A(B[2]), .ZN(n280) );
  NAND2_X1 U277 ( .A1(B[2]), .A2(n274), .ZN(n77) );
  XNOR2_X1 U278 ( .A(n50), .B(n51), .ZN(DIFF[8]) );
  INV_X1 U279 ( .A(n64), .ZN(n62) );
  INV_X1 U280 ( .A(n65), .ZN(n61) );
  XNOR2_X1 U281 ( .A(n67), .B(n65), .ZN(DIFF[5]) );
  INV_X1 U282 ( .A(n71), .ZN(n68) );
  OAI21_X1 U283 ( .B1(n75), .B2(n76), .A(n4), .ZN(n74) );
  INV_X1 U284 ( .A(n77), .ZN(n76) );
  INV_X1 U285 ( .A(n78), .ZN(n75) );
  INV_X1 U286 ( .A(n91), .ZN(n89) );
  INV_X1 U287 ( .A(n94), .ZN(n93) );
  INV_X1 U288 ( .A(net15475), .ZN(net15471) );
  NAND3_X1 U289 ( .A1(n91), .A2(n86), .A3(n92), .ZN(net15462) );
  NOR2_X1 U290 ( .A1(n97), .A2(n45), .ZN(n96) );
  INV_X1 U291 ( .A(n86), .ZN(n97) );
  INV_X1 U292 ( .A(n90), .ZN(n101) );
  INV_X1 U293 ( .A(n116), .ZN(n115) );
  INV_X1 U294 ( .A(n123), .ZN(n122) );
  INV_X1 U295 ( .A(n124), .ZN(n120) );
  NAND3_X1 U296 ( .A1(n125), .A2(n113), .A3(n121), .ZN(net15500) );
  XNOR2_X1 U297 ( .A(n126), .B(n127), .ZN(DIFF[23]) );
  INV_X1 U298 ( .A(n125), .ZN(n118) );
  XNOR2_X1 U299 ( .A(n141), .B(n38), .ZN(DIFF[20]) );
  INV_X1 U300 ( .A(n148), .ZN(n147) );
  INV_X1 U301 ( .A(n155), .ZN(n154) );
  INV_X1 U302 ( .A(n156), .ZN(n152) );
  NAND3_X1 U303 ( .A1(n157), .A2(n145), .A3(n153), .ZN(n143) );
  XNOR2_X1 U304 ( .A(n163), .B(n164), .ZN(DIFF[19]) );
  OAI21_X1 U305 ( .B1(n165), .B2(n150), .A(n151), .ZN(n164) );
  INV_X1 U306 ( .A(n157), .ZN(n150) );
  INV_X1 U307 ( .A(n166), .ZN(n165) );
  XNOR2_X1 U308 ( .A(n179), .B(n41), .ZN(DIFF[16]) );
  NAND4_X1 U309 ( .A1(n2), .A2(n184), .A3(n185), .A4(n33), .ZN(n183) );
  INV_X1 U310 ( .A(n186), .ZN(n185) );
  INV_X1 U311 ( .A(n191), .ZN(n190) );
  INV_X1 U312 ( .A(n198), .ZN(n197) );
  INV_X1 U313 ( .A(n199), .ZN(n195) );
  NAND3_X1 U314 ( .A1(n200), .A2(n33), .A3(n201), .ZN(n181) );
  INV_X1 U315 ( .A(n202), .ZN(n184) );
  INV_X1 U316 ( .A(n208), .ZN(n193) );
  INV_X1 U317 ( .A(n214), .ZN(n213) );
  INV_X1 U318 ( .A(n196), .ZN(n219) );
  INV_X1 U319 ( .A(n220), .ZN(n218) );
  XNOR2_X1 U320 ( .A(n223), .B(n220), .ZN(DIFF[13]) );
  INV_X1 U321 ( .A(n226), .ZN(n225) );
  INV_X1 U322 ( .A(n207), .ZN(n224) );
  INV_X1 U323 ( .A(n204), .ZN(n230) );
  INV_X1 U324 ( .A(n237), .ZN(n236) );
  INV_X1 U325 ( .A(n238), .ZN(n234) );
  INV_X1 U326 ( .A(n51), .ZN(n229) );
  XNOR2_X1 U327 ( .A(n243), .B(n244), .ZN(DIFF[11]) );
  INV_X1 U328 ( .A(n239), .ZN(n246) );
  INV_X1 U329 ( .A(n247), .ZN(n245) );
  XNOR2_X1 U330 ( .A(n250), .B(n247), .ZN(DIFF[10]) );
  INV_X1 U331 ( .A(n27), .ZN(n256) );
  INV_X1 U332 ( .A(n57), .ZN(n262) );
  INV_X1 U333 ( .A(n73), .ZN(n69) );
  NAND3_X1 U334 ( .A1(n79), .A2(n77), .A3(n269), .ZN(n186) );
  NOR2_X1 U335 ( .A1(n270), .A2(n36), .ZN(n269) );
  INV_X1 U336 ( .A(n84), .ZN(n270) );
  INV_X1 U337 ( .A(n80), .ZN(n277) );
  INV_X1 U338 ( .A(n48), .ZN(n251) );
endmodule


module ALU_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240;

  INV_X1 U2 ( .A(n86), .ZN(n19) );
  INV_X1 U3 ( .A(n16), .ZN(n202) );
  OAI21_X1 U4 ( .B1(n232), .B2(n181), .A(n227), .ZN(n41) );
  INV_X1 U5 ( .A(n13), .ZN(n181) );
  CLKBUF_X1 U6 ( .A(n77), .Z(n21) );
  NAND2_X1 U7 ( .A1(B[6]), .A2(A[6]), .ZN(n1) );
  OR2_X1 U8 ( .A1(B[5]), .A2(A[5]), .ZN(n2) );
  OR2_X1 U9 ( .A1(B[6]), .A2(A[6]), .ZN(n3) );
  NAND2_X1 U10 ( .A1(B[4]), .A2(A[4]), .ZN(n4) );
  NAND2_X1 U11 ( .A1(B[5]), .A2(A[5]), .ZN(n5) );
  BUF_X1 U12 ( .A(n43), .Z(n6) );
  OR2_X1 U13 ( .A1(B[14]), .A2(A[14]), .ZN(n7) );
  AND2_X1 U14 ( .A1(B[6]), .A2(A[6]), .ZN(n8) );
  CLKBUF_X1 U15 ( .A(n177), .Z(n9) );
  NAND2_X1 U16 ( .A1(B[1]), .A2(A[1]), .ZN(n10) );
  NAND2_X1 U17 ( .A1(B[8]), .A2(A[8]), .ZN(n11) );
  CLKBUF_X1 U18 ( .A(n47), .Z(n12) );
  AND4_X2 U19 ( .A1(n3), .A2(n2), .A3(n60), .A4(n49), .ZN(n13) );
  CLKBUF_X1 U20 ( .A(n216), .Z(n14) );
  OR2_X1 U21 ( .A1(B[10]), .A2(A[10]), .ZN(n216) );
  CLKBUF_X1 U22 ( .A(n157), .Z(n15) );
  OR2_X2 U23 ( .A1(B[11]), .A2(A[11]), .ZN(n214) );
  AND2_X1 U24 ( .A1(n204), .A2(n196), .ZN(n16) );
  CLKBUF_X1 U25 ( .A(n90), .Z(n17) );
  CLKBUF_X1 U26 ( .A(n140), .Z(n18) );
  NOR2_X1 U27 ( .A1(n20), .A2(n19), .ZN(n77) );
  AND2_X1 U28 ( .A1(n28), .A2(n88), .ZN(n20) );
  CLKBUF_X1 U29 ( .A(n180), .Z(n22) );
  CLKBUF_X1 U30 ( .A(B[0]), .Z(n23) );
  OAI21_X1 U31 ( .B1(n18), .B2(n141), .A(n142), .ZN(n24) );
  OAI21_X1 U32 ( .B1(n140), .B2(n141), .A(n142), .ZN(n137) );
  CLKBUF_X1 U33 ( .A(n115), .Z(n25) );
  CLKBUF_X1 U34 ( .A(n167), .Z(n26) );
  OAI21_X1 U35 ( .B1(n115), .B2(n116), .A(n117), .ZN(n27) );
  OAI21_X1 U36 ( .B1(n90), .B2(n91), .A(n92), .ZN(n28) );
  OAI21_X1 U37 ( .B1(n76), .B2(n21), .A(n78), .ZN(n29) );
  XOR2_X1 U38 ( .A(n30), .B(n21), .Z(SUM[29]) );
  NAND2_X1 U39 ( .A1(n78), .A2(n79), .ZN(n30) );
  XOR2_X1 U40 ( .A(B[31]), .B(A[31]), .Z(n31) );
  OR2_X1 U41 ( .A1(B[2]), .A2(A[2]), .ZN(n85) );
  AND2_X1 U42 ( .A1(n15), .A2(n233), .ZN(SUM[0]) );
  OAI21_X1 U43 ( .B1(n207), .B2(n9), .A(n208), .ZN(n205) );
  AOI22_X1 U44 ( .A1(n173), .A2(n174), .B1(n176), .B2(n175), .ZN(n172) );
  NOR2_X1 U45 ( .A1(n186), .A2(n187), .ZN(n170) );
  NAND4_X1 U46 ( .A1(n180), .A2(n175), .A3(n13), .A4(n179), .ZN(n171) );
  INV_X1 U47 ( .A(n23), .ZN(n239) );
  NOR2_X1 U48 ( .A1(n177), .A2(n178), .ZN(n173) );
  XNOR2_X1 U49 ( .A(n114), .B(n33), .ZN(SUM[24]) );
  XNOR2_X1 U50 ( .A(n206), .B(n205), .ZN(SUM[12]) );
  XNOR2_X1 U51 ( .A(n111), .B(n110), .ZN(SUM[25]) );
  XNOR2_X1 U52 ( .A(n203), .B(n202), .ZN(SUM[13]) );
  XNOR2_X1 U53 ( .A(n201), .B(n200), .ZN(SUM[14]) );
  XNOR2_X1 U54 ( .A(n106), .B(n108), .ZN(SUM[26]) );
  XNOR2_X1 U55 ( .A(n166), .B(n165), .ZN(SUM[17]) );
  XNOR2_X1 U56 ( .A(n163), .B(n162), .ZN(SUM[18]) );
  XNOR2_X1 U57 ( .A(n136), .B(n135), .ZN(SUM[21]) );
  XNOR2_X1 U58 ( .A(n131), .B(n133), .ZN(SUM[22]) );
  OAI21_X1 U59 ( .B1(n16), .B2(n195), .A(n194), .ZN(n200) );
  OAI21_X1 U60 ( .B1(n52), .B2(n53), .A(n5), .ZN(n48) );
  OAI21_X1 U61 ( .B1(n224), .B2(n225), .A(n39), .ZN(n222) );
  NAND4_X1 U62 ( .A1(n216), .A2(n214), .A3(n38), .A4(n43), .ZN(n177) );
  OAI211_X1 U63 ( .C1(n209), .C2(n210), .A(n211), .B(n212), .ZN(n176) );
  NAND2_X1 U64 ( .A1(n213), .A2(n214), .ZN(n211) );
  NAND2_X1 U65 ( .A1(n214), .A2(n38), .ZN(n210) );
  NAND2_X1 U66 ( .A1(n216), .A2(n217), .ZN(n209) );
  NOR2_X1 U67 ( .A1(n143), .A2(n144), .ZN(n142) );
  NAND2_X1 U68 ( .A1(n212), .A2(n214), .ZN(n218) );
  NAND2_X1 U69 ( .A1(n68), .A2(n69), .ZN(n62) );
  AOI21_X1 U70 ( .B1(n122), .B2(n131), .A(n132), .ZN(n129) );
  OAI21_X1 U71 ( .B1(n17), .B2(n91), .A(n92), .ZN(n87) );
  NOR2_X1 U72 ( .A1(n34), .A2(n93), .ZN(n92) );
  AOI21_X1 U73 ( .B1(n94), .B2(n95), .A(n96), .ZN(n93) );
  OAI21_X1 U74 ( .B1(n25), .B2(n116), .A(n117), .ZN(n112) );
  NOR2_X1 U75 ( .A1(n35), .A2(n118), .ZN(n117) );
  AOI21_X1 U76 ( .B1(n119), .B2(n120), .A(n121), .ZN(n118) );
  AOI21_X1 U77 ( .B1(n189), .B2(n190), .A(n191), .ZN(n186) );
  OAI21_X1 U78 ( .B1(n192), .B2(n193), .A(n7), .ZN(n189) );
  INV_X1 U79 ( .A(n194), .ZN(n193) );
  XNOR2_X1 U80 ( .A(n129), .B(n130), .ZN(SUM[23]) );
  NAND4_X1 U81 ( .A1(n182), .A2(n183), .A3(n184), .A4(n185), .ZN(n178) );
  AOI21_X1 U82 ( .B1(n145), .B2(n146), .A(n147), .ZN(n144) );
  NAND2_X1 U83 ( .A1(n149), .A2(n150), .ZN(n145) );
  OAI21_X1 U84 ( .B1(n151), .B2(n152), .A(n153), .ZN(n150) );
  OAI21_X1 U85 ( .B1(n77), .B2(n76), .A(n78), .ZN(n71) );
  NOR2_X1 U86 ( .A1(n121), .A2(n35), .ZN(n130) );
  NAND2_X1 U87 ( .A1(n228), .A2(n229), .ZN(n174) );
  AOI21_X1 U88 ( .B1(n8), .B2(n49), .A(n231), .ZN(n228) );
  NAND4_X1 U89 ( .A1(n230), .A2(n55), .A3(n47), .A4(n49), .ZN(n229) );
  NAND2_X1 U90 ( .A1(n25), .A2(n125), .ZN(n135) );
  NAND2_X1 U91 ( .A1(n18), .A2(n152), .ZN(n165) );
  NAND2_X1 U92 ( .A1(n235), .A2(n234), .ZN(n180) );
  AOI21_X1 U93 ( .B1(n237), .B2(n68), .A(n238), .ZN(n234) );
  NAND4_X1 U94 ( .A1(n236), .A2(n83), .A3(n85), .A4(n68), .ZN(n235) );
  NAND2_X1 U95 ( .A1(n58), .A2(n4), .ZN(n56) );
  NAND2_X1 U96 ( .A1(n22), .A2(n60), .ZN(n58) );
  XNOR2_X1 U97 ( .A(n61), .B(n22), .ZN(SUM[4]) );
  NOR2_X1 U98 ( .A1(n195), .A2(n196), .ZN(n192) );
  NAND2_X1 U99 ( .A1(n134), .A2(n126), .ZN(n131) );
  NAND2_X1 U100 ( .A1(n127), .A2(n135), .ZN(n134) );
  NAND2_X1 U101 ( .A1(n17), .A2(n100), .ZN(n110) );
  NAND2_X1 U102 ( .A1(n109), .A2(n101), .ZN(n106) );
  NAND2_X1 U103 ( .A1(n102), .A2(n110), .ZN(n109) );
  NAND2_X1 U104 ( .A1(n226), .A2(n11), .ZN(n37) );
  NAND2_X1 U105 ( .A1(n41), .A2(n6), .ZN(n226) );
  NAND2_X1 U106 ( .A1(n205), .A2(n182), .ZN(n204) );
  NAND2_X1 U107 ( .A1(n164), .A2(n153), .ZN(n162) );
  NAND2_X1 U108 ( .A1(n154), .A2(n165), .ZN(n164) );
  XNOR2_X1 U109 ( .A(n104), .B(n105), .ZN(SUM[27]) );
  NOR2_X1 U110 ( .A1(n96), .A2(n34), .ZN(n105) );
  AOI21_X1 U111 ( .B1(n97), .B2(n106), .A(n107), .ZN(n104) );
  INV_X1 U112 ( .A(n15), .ZN(n84) );
  XNOR2_X1 U113 ( .A(n44), .B(n45), .ZN(SUM[7]) );
  NAND2_X1 U114 ( .A1(n49), .A2(n50), .ZN(n44) );
  NAND2_X1 U115 ( .A1(n46), .A2(n1), .ZN(n45) );
  NAND2_X1 U116 ( .A1(n12), .A2(n48), .ZN(n46) );
  XNOR2_X1 U117 ( .A(n40), .B(n41), .ZN(SUM[8]) );
  NAND2_X1 U118 ( .A1(n11), .A2(n6), .ZN(n40) );
  XNOR2_X1 U119 ( .A(n51), .B(n48), .ZN(SUM[6]) );
  NAND2_X1 U120 ( .A1(n12), .A2(n1), .ZN(n51) );
  XNOR2_X1 U121 ( .A(n36), .B(n37), .ZN(SUM[9]) );
  NAND2_X1 U122 ( .A1(n38), .A2(n39), .ZN(n36) );
  XNOR2_X1 U123 ( .A(n223), .B(n222), .ZN(SUM[10]) );
  NAND2_X1 U124 ( .A1(n215), .A2(n14), .ZN(n223) );
  XNOR2_X1 U125 ( .A(n57), .B(n56), .ZN(SUM[5]) );
  NAND2_X1 U126 ( .A1(n2), .A2(n5), .ZN(n57) );
  XNOR2_X1 U127 ( .A(n87), .B(n89), .ZN(SUM[28]) );
  NAND2_X1 U128 ( .A1(n86), .A2(n88), .ZN(n89) );
  XNOR2_X1 U129 ( .A(n80), .B(n67), .ZN(SUM[2]) );
  NAND2_X1 U130 ( .A1(n85), .A2(n66), .ZN(n80) );
  XNOR2_X1 U131 ( .A(n29), .B(n75), .ZN(SUM[30]) );
  NAND2_X1 U132 ( .A1(n74), .A2(n72), .ZN(n75) );
  NAND2_X1 U133 ( .A1(n167), .A2(n168), .ZN(n140) );
  NAND2_X1 U134 ( .A1(n4), .A2(n60), .ZN(n61) );
  NAND2_X1 U135 ( .A1(n137), .A2(n138), .ZN(n115) );
  NAND2_X1 U136 ( .A1(n27), .A2(n113), .ZN(n90) );
  NAND2_X1 U137 ( .A1(n54), .A2(n59), .ZN(n230) );
  XNOR2_X1 U138 ( .A(n197), .B(n198), .ZN(SUM[15]) );
  NAND2_X1 U139 ( .A1(n188), .A2(n185), .ZN(n197) );
  NAND2_X1 U140 ( .A1(n190), .A2(n199), .ZN(n198) );
  NAND2_X1 U141 ( .A1(n7), .A2(n200), .ZN(n199) );
  NAND2_X1 U142 ( .A1(n39), .A2(n42), .ZN(n217) );
  NAND2_X1 U143 ( .A1(n95), .A2(n97), .ZN(n108) );
  NAND2_X1 U144 ( .A1(n120), .A2(n122), .ZN(n133) );
  NAND2_X1 U145 ( .A1(n196), .A2(n182), .ZN(n206) );
  NAND2_X1 U146 ( .A1(n153), .A2(n154), .ZN(n166) );
  NAND2_X1 U147 ( .A1(n190), .A2(n7), .ZN(n201) );
  NAND2_X1 U148 ( .A1(n194), .A2(n183), .ZN(n203) );
  NAND2_X1 U149 ( .A1(n157), .A2(n82), .ZN(n236) );
  NAND2_X1 U150 ( .A1(n126), .A2(n127), .ZN(n136) );
  NAND2_X1 U151 ( .A1(n83), .A2(n10), .ZN(n156) );
  NAND2_X1 U152 ( .A1(n146), .A2(n149), .ZN(n163) );
  NAND2_X1 U153 ( .A1(n101), .A2(n102), .ZN(n111) );
  NAND2_X1 U154 ( .A1(n125), .A2(n138), .ZN(n139) );
  NAND2_X1 U155 ( .A1(n152), .A2(n168), .ZN(n169) );
  NAND2_X1 U156 ( .A1(n122), .A2(n123), .ZN(n119) );
  OAI21_X1 U157 ( .B1(n124), .B2(n125), .A(n126), .ZN(n123) );
  INV_X1 U158 ( .A(n188), .ZN(n187) );
  NAND2_X1 U159 ( .A1(n97), .A2(n98), .ZN(n94) );
  OAI21_X1 U160 ( .B1(n99), .B2(n100), .A(n101), .ZN(n98) );
  NAND2_X1 U161 ( .A1(n81), .A2(n10), .ZN(n67) );
  NAND2_X1 U162 ( .A1(n83), .A2(n84), .ZN(n81) );
  NAND2_X1 U163 ( .A1(n155), .A2(n148), .ZN(n158) );
  AND2_X1 U164 ( .A1(n100), .A2(n113), .ZN(n33) );
  NAND2_X1 U165 ( .A1(B[0]), .A2(A[0]), .ZN(n157) );
  NAND2_X1 U166 ( .A1(B[5]), .A2(A[5]), .ZN(n54) );
  NAND2_X1 U167 ( .A1(B[8]), .A2(A[8]), .ZN(n42) );
  NAND2_X1 U168 ( .A1(B[20]), .A2(A[20]), .ZN(n125) );
  NAND2_X1 U169 ( .A1(B[9]), .A2(A[9]), .ZN(n39) );
  NAND2_X1 U170 ( .A1(B[12]), .A2(A[12]), .ZN(n196) );
  NAND2_X1 U171 ( .A1(B[16]), .A2(A[16]), .ZN(n152) );
  NAND2_X1 U172 ( .A1(B[17]), .A2(A[17]), .ZN(n153) );
  NAND2_X1 U173 ( .A1(B[30]), .A2(A[30]), .ZN(n74) );
  NAND2_X1 U174 ( .A1(B[14]), .A2(A[14]), .ZN(n190) );
  NAND2_X1 U175 ( .A1(B[13]), .A2(A[13]), .ZN(n194) );
  OR2_X1 U176 ( .A1(B[7]), .A2(A[7]), .ZN(n49) );
  NAND2_X1 U177 ( .A1(B[21]), .A2(A[21]), .ZN(n126) );
  NAND2_X1 U178 ( .A1(B[10]), .A2(A[10]), .ZN(n215) );
  NAND2_X1 U179 ( .A1(B[18]), .A2(A[18]), .ZN(n146) );
  NAND2_X1 U180 ( .A1(B[25]), .A2(A[25]), .ZN(n101) );
  NAND2_X1 U181 ( .A1(B[26]), .A2(A[26]), .ZN(n95) );
  NAND2_X1 U182 ( .A1(B[11]), .A2(A[11]), .ZN(n212) );
  OR2_X1 U183 ( .A1(B[14]), .A2(A[14]), .ZN(n184) );
  NAND2_X1 U184 ( .A1(B[22]), .A2(A[22]), .ZN(n120) );
  NAND2_X1 U185 ( .A1(B[1]), .A2(A[1]), .ZN(n82) );
  NAND2_X1 U186 ( .A1(B[15]), .A2(A[15]), .ZN(n188) );
  OR2_X1 U187 ( .A1(B[9]), .A2(A[9]), .ZN(n38) );
  NAND2_X1 U188 ( .A1(B[7]), .A2(A[7]), .ZN(n50) );
  NAND2_X1 U189 ( .A1(B[24]), .A2(A[24]), .ZN(n100) );
  OR2_X1 U190 ( .A1(B[26]), .A2(A[26]), .ZN(n97) );
  NAND2_X1 U191 ( .A1(B[3]), .A2(A[3]), .ZN(n69) );
  NAND2_X1 U192 ( .A1(B[19]), .A2(A[19]), .ZN(n155) );
  AND2_X1 U193 ( .A1(B[27]), .A2(A[27]), .ZN(n34) );
  AND2_X1 U194 ( .A1(B[23]), .A2(A[23]), .ZN(n35) );
  OR2_X1 U195 ( .A1(B[3]), .A2(A[3]), .ZN(n68) );
  OR2_X1 U196 ( .A1(B[25]), .A2(A[25]), .ZN(n102) );
  OR2_X1 U197 ( .A1(B[17]), .A2(A[17]), .ZN(n154) );
  OR2_X1 U198 ( .A1(B[18]), .A2(A[18]), .ZN(n149) );
  NAND2_X1 U199 ( .A1(B[28]), .A2(A[28]), .ZN(n86) );
  OR2_X1 U200 ( .A1(B[12]), .A2(A[12]), .ZN(n182) );
  OR2_X1 U201 ( .A1(B[4]), .A2(A[4]), .ZN(n60) );
  OR2_X1 U202 ( .A1(B[30]), .A2(A[30]), .ZN(n72) );
  NAND2_X1 U203 ( .A1(B[29]), .A2(A[29]), .ZN(n78) );
  XNOR2_X1 U204 ( .A(n156), .B(n84), .ZN(SUM[1]) );
  OR2_X1 U205 ( .A1(B[13]), .A2(A[13]), .ZN(n183) );
  XNOR2_X1 U206 ( .A(n70), .B(n31), .ZN(SUM[31]) );
  OR2_X1 U207 ( .A1(B[5]), .A2(A[5]), .ZN(n55) );
  OR2_X1 U208 ( .A1(B[19]), .A2(A[19]), .ZN(n148) );
  OR2_X1 U209 ( .A1(B[20]), .A2(A[20]), .ZN(n138) );
  OR2_X1 U210 ( .A1(B[28]), .A2(A[28]), .ZN(n88) );
  OR2_X1 U211 ( .A1(B[6]), .A2(A[6]), .ZN(n47) );
  OR2_X1 U212 ( .A1(B[8]), .A2(A[8]), .ZN(n43) );
  OR2_X1 U213 ( .A1(B[16]), .A2(A[16]), .ZN(n168) );
  OR2_X1 U214 ( .A1(B[15]), .A2(A[15]), .ZN(n185) );
  OR2_X1 U215 ( .A1(B[27]), .A2(A[27]), .ZN(n103) );
  OR2_X1 U216 ( .A1(B[23]), .A2(A[23]), .ZN(n128) );
  OR2_X1 U217 ( .A1(B[1]), .A2(A[1]), .ZN(n83) );
  OR2_X1 U218 ( .A1(B[24]), .A2(A[24]), .ZN(n113) );
  OR2_X1 U219 ( .A1(B[29]), .A2(A[29]), .ZN(n79) );
  OR2_X1 U220 ( .A1(B[21]), .A2(A[21]), .ZN(n127) );
  OR2_X1 U221 ( .A1(B[22]), .A2(A[22]), .ZN(n122) );
  NAND2_X1 U222 ( .A1(n239), .A2(n240), .ZN(n233) );
  INV_X1 U223 ( .A(A[0]), .ZN(n240) );
  NAND3_X1 U224 ( .A1(n171), .A2(n170), .A3(n172), .ZN(n167) );
  NAND2_X1 U225 ( .A1(B[2]), .A2(A[2]), .ZN(n66) );
  NAND2_X1 U226 ( .A1(B[4]), .A2(A[4]), .ZN(n59) );
  INV_X1 U227 ( .A(n2), .ZN(n53) );
  INV_X1 U228 ( .A(n56), .ZN(n52) );
  XNOR2_X1 U229 ( .A(n62), .B(n63), .ZN(SUM[3]) );
  OAI21_X1 U230 ( .B1(n64), .B2(n65), .A(n66), .ZN(n63) );
  INV_X1 U231 ( .A(n67), .ZN(n64) );
  AOI21_X1 U232 ( .B1(n71), .B2(n72), .A(n73), .ZN(n70) );
  INV_X1 U233 ( .A(n74), .ZN(n73) );
  INV_X1 U234 ( .A(n79), .ZN(n76) );
  INV_X1 U235 ( .A(n102), .ZN(n99) );
  NAND3_X1 U236 ( .A1(n97), .A2(n103), .A3(n102), .ZN(n91) );
  INV_X1 U237 ( .A(n103), .ZN(n96) );
  INV_X1 U238 ( .A(n95), .ZN(n107) );
  INV_X1 U239 ( .A(n112), .ZN(n114) );
  INV_X1 U240 ( .A(n127), .ZN(n124) );
  NAND3_X1 U241 ( .A1(n122), .A2(n128), .A3(n127), .ZN(n116) );
  INV_X1 U242 ( .A(n128), .ZN(n121) );
  INV_X1 U243 ( .A(n120), .ZN(n132) );
  XNOR2_X1 U244 ( .A(n139), .B(n24), .ZN(SUM[20]) );
  INV_X1 U245 ( .A(n148), .ZN(n147) );
  INV_X1 U246 ( .A(n154), .ZN(n151) );
  INV_X1 U247 ( .A(n155), .ZN(n143) );
  NAND3_X1 U248 ( .A1(n149), .A2(n148), .A3(n154), .ZN(n141) );
  XNOR2_X1 U249 ( .A(n158), .B(n159), .ZN(SUM[19]) );
  OAI21_X1 U250 ( .B1(n160), .B2(n161), .A(n146), .ZN(n159) );
  INV_X1 U251 ( .A(n149), .ZN(n161) );
  INV_X1 U252 ( .A(n162), .ZN(n160) );
  XNOR2_X1 U253 ( .A(n169), .B(n26), .ZN(SUM[16]) );
  INV_X1 U254 ( .A(n178), .ZN(n175) );
  INV_X1 U255 ( .A(n177), .ZN(n179) );
  INV_X1 U256 ( .A(n185), .ZN(n191) );
  INV_X1 U257 ( .A(n183), .ZN(n195) );
  INV_X1 U258 ( .A(n176), .ZN(n208) );
  INV_X1 U259 ( .A(n215), .ZN(n213) );
  INV_X1 U260 ( .A(n41), .ZN(n207) );
  XNOR2_X1 U261 ( .A(n218), .B(n219), .ZN(SUM[11]) );
  OAI21_X1 U262 ( .B1(n220), .B2(n221), .A(n215), .ZN(n219) );
  INV_X1 U263 ( .A(n14), .ZN(n221) );
  INV_X1 U264 ( .A(n222), .ZN(n220) );
  INV_X1 U265 ( .A(n37), .ZN(n225) );
  INV_X1 U266 ( .A(n174), .ZN(n227) );
  INV_X1 U267 ( .A(n50), .ZN(n231) );
  INV_X1 U268 ( .A(n85), .ZN(n65) );
  INV_X1 U269 ( .A(n22), .ZN(n232) );
  INV_X1 U270 ( .A(n69), .ZN(n238) );
  INV_X1 U271 ( .A(n66), .ZN(n237) );
  INV_X1 U272 ( .A(n38), .ZN(n224) );
endmodule


module ALU ( OP1, OP2, ALU_OP, RES, ZERO );
  input [31:0] OP1;
  input [31:0] OP2;
  input [3:0] ALU_OP;
  output [31:0] RES;
  output ZERO;
  wire   N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N189, N191,
         N193, n124, n125, n126, n127, n128, n142, n143, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n205, n206, n207, n208, n209, n210, n211, n212, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n231, n232, n234, n235,
         n236, n237, n238, n239, n240, n242, n243, n244, n245, n252, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n271, n272,
         n273, n274, n275, n276, n277, n278, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n298, n299, n300, n301, n302, n303, n304,
         n305, n312, n313, n314, n315, n316, n317, n318, n319, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n344, n345, n346, n347, n348, n349, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n386, n387, n388, n389, n390, n391, n392, n393, n400,
         n401, n402, n403, n404, n405, n406, n407, n414, n415, n416, n423,
         n424, n425, n426, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n446, n447, n448, n449, n456, n457, n458, n459, n460, n467,
         n468, n469, n470, n477, n478, n479, n480, n487, n488, n489, n490,
         n491, n498, n499, n500, n501, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n524, n525, n526, n527, n528, n529, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n565, n573, n574, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n144, n159, n160, n161, n162, n174, n175, n176, n188, n189, n190,
         n202, n203, n204, n213, n214, n215, n226, n227, n228, n229, n230,
         n233, n241, n246, n247, n248, n249, n250, n251, n253, n254, n265,
         n266, n267, n268, n269, n270, n279, n280, n281, n282, n292, n293,
         n294, n295, n296, n297, n306, n307, n308, n309, n310, n311, n320,
         n321, n322, n323, n324, n338, n339, n340, n341, n342, n343, n350,
         n351, n352, n353, n354, n355, n365, n366, n367, n368, n369, n370,
         n380, n381, n382, n383, n384, n385, n394, n395, n396, n397, n398,
         n399, n408, n409, n410, n411, n412, n413, n417, n418, n419, n420,
         n421, n422, n427, n428, n429, n430, n431, n441, n442, n443, n444,
         n445, n450, n451, n452, n453, n454, n455, n461, n462, n463, n464,
         n465, n466, n471, n472, n473, n474, n475, n476, n481, n482, n483,
         n484, n485, n486, n492, n493, n494, n495, n496, n497, n502, n503,
         n504, n505, n506, n507, n518, n519, n520, n521, n522, n523, n530,
         n531, n532, n533, n548, n549, n550, n563, n564, n566, n567, n568,
         n569, n570, n571, n572, n575, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711;

  NAND2_X2 U432 ( .A1(n710), .A2(n697), .ZN(n331) );
  NAND2_X2 U442 ( .A1(n6), .A2(n697), .ZN(n147) );
  OAI33_X1 U626 ( .A1(n100), .A2(n18), .A3(n709), .B1(n578), .B2(n579), .B3(
        n235), .ZN(n577) );
  NAND3_X1 U627 ( .A1(n73), .A2(n51), .A3(n698), .ZN(n592) );
  ALU_DW01_cmp6_0 r131 ( .A(OP1), .B({OP2[31:2], n16, OP2[0]}), .TC(1'b0), 
        .LE(N189), .GE(N191), .NE(N193) );
  ALU_DW01_sub_2 sub_30 ( .A(OP1), .B({OP2[31:27], n15, OP2[25:23], n14, 
        OP2[21], n33, OP2[19:3], n38, OP2[1:0]}), .CI(1'b0), .DIFF({N187, N186, 
        N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, 
        N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, 
        N161, N160, N159, N158, N157, N156}) );
  ALU_DW01_add_2 add_28 ( .A({OP1[31:2], n45, n18}), .B({OP2[31:27], n15, 
        OP2[25:23], n14, OP2[21], n33, OP2[19:15], n24, OP2[13:9], n23, 
        OP2[7:6], n22, n30, OP2[3], n38, n16, n63}), .CI(1'b0), .SUM({N154, 
        N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, 
        N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, 
        N129, N128, N127, N126, N125, N124, N123}) );
  OAI221_X4 U6 ( .B1(n92), .B2(n618), .C1(n91), .C2(n619), .A(n588), .ZN(n378)
         );
  OAI221_X1 U7 ( .B1(n89), .B2(n693), .C1(n257), .C2(n695), .A(n582), .ZN(n581) );
  OAI221_X1 U8 ( .B1(n94), .B2(n621), .C1(n91), .C2(n622), .A(n510), .ZN(n364)
         );
  OAI221_X1 U9 ( .B1(n93), .B2(n696), .C1(n91), .C2(n695), .A(n546), .ZN(n237)
         );
  OAI221_X1 U10 ( .B1(n94), .B2(n636), .C1(n91), .C2(n637), .A(n558), .ZN(n196) );
  OAI221_X1 U11 ( .B1(n94), .B2(n632), .C1(n91), .C2(n633), .A(n557), .ZN(n198) );
  OAI221_X1 U12 ( .B1(n94), .B2(n637), .C1(n91), .C2(n674), .A(n439), .ZN(n156) );
  OAI221_X1 U13 ( .B1(n94), .B2(n635), .C1(n91), .C2(n634), .A(n469), .ZN(n303) );
  OAI221_X1 U14 ( .B1(n95), .B2(n632), .C1(n91), .C2(n631), .A(n426), .ZN(n316) );
  OAI221_X1 U15 ( .B1(n92), .B2(n674), .C1(n91), .C2(n637), .A(n501), .ZN(n347) );
  OAI221_X1 U16 ( .B1(n94), .B2(n682), .C1(n91), .C2(n680), .A(n561), .ZN(n402) );
  OAI221_X1 U17 ( .B1(n94), .B2(n690), .C1(n91), .C2(n688), .A(n560), .ZN(n404) );
  AOI221_X1 U18 ( .B1(n407), .B2(n705), .C1(n406), .C2(n74), .A(n459), .ZN(
        n291) );
  OAI221_X1 U19 ( .B1(n92), .B2(n630), .C1(n91), .C2(n631), .A(n589), .ZN(n170) );
  OAI221_X1 U20 ( .B1(n92), .B2(n634), .C1(n91), .C2(n635), .A(n585), .ZN(n168) );
  OAI221_X1 U21 ( .B1(n94), .B2(n674), .C1(n91), .C2(n676), .A(n586), .ZN(n171) );
  OAI221_X1 U22 ( .B1(n89), .B2(n620), .C1(n257), .C2(n619), .A(n258), .ZN(
        n256) );
  AOI211_X1 U23 ( .C1(n47), .C2(n57), .A(n225), .B(n215), .ZN(n121) );
  AOI211_X1 U24 ( .C1(n2), .C2(n57), .A(n201), .B(n215), .ZN(n134) );
  AOI211_X1 U25 ( .C1(OP2[10]), .C2(n57), .A(n562), .B(n215), .ZN(n188) );
  AOI221_X1 U26 ( .B1(n379), .B2(n705), .C1(n169), .C2(n74), .A(n3), .ZN(n26)
         );
  AOI211_X1 U27 ( .C1(n32), .C2(n57), .A(n173), .B(n215), .ZN(n144) );
  INV_X1 U28 ( .A(OP2[6]), .ZN(n1) );
  INV_X1 U29 ( .A(n1), .ZN(n2) );
  CLKBUF_X1 U30 ( .A(n587), .Z(n3) );
  CLKBUF_X1 U31 ( .A(n42), .Z(n4) );
  INV_X2 U32 ( .A(n58), .ZN(n90) );
  OAI221_X1 U33 ( .B1(n92), .B2(n637), .C1(n90), .C2(n636), .A(n491), .ZN(n329) );
  OAI221_X1 U34 ( .B1(n93), .B2(n678), .C1(n90), .C2(n676), .A(n528), .ZN(n373) );
  OAI221_X4 U35 ( .B1(n94), .B2(n633), .C1(n91), .C2(n632), .A(n449), .ZN(n263) );
  OAI221_X4 U36 ( .B1(n93), .B2(n680), .C1(n91), .C2(n678), .A(n545), .ZN(n387) );
  OAI221_X4 U37 ( .B1(n93), .B2(n688), .C1(n91), .C2(n686), .A(n544), .ZN(n391) );
  OAI221_X4 U38 ( .B1(n94), .B2(n620), .C1(n91), .C2(n621), .A(n559), .ZN(n407) );
  OAI221_X4 U39 ( .B1(n92), .B2(n628), .C1(n91), .C2(n629), .A(n555), .ZN(n197) );
  OAI221_X1 U40 ( .B1(n94), .B2(n676), .C1(n90), .C2(n674), .A(n515), .ZN(n358) );
  OAI221_X1 U41 ( .B1(n92), .B2(n629), .C1(n90), .C2(n630), .A(n513), .ZN(n155) );
  INV_X2 U42 ( .A(n58), .ZN(n89) );
  AND2_X1 U43 ( .A1(OP1[31]), .A2(n82), .ZN(n5) );
  AND2_X1 U44 ( .A1(n593), .A2(n574), .ZN(n6) );
  BUF_X1 U45 ( .A(OP1[0]), .Z(n18) );
  AND2_X1 U46 ( .A1(n593), .A2(n62), .ZN(n7) );
  AND3_X1 U47 ( .A1(n580), .A2(n638), .A3(ALU_OP[0]), .ZN(n8) );
  NAND2_X1 U48 ( .A1(N156), .A2(n68), .ZN(n9) );
  CLKBUF_X1 U49 ( .A(OP2[13]), .Z(n10) );
  BUF_X2 U50 ( .A(OP2[4]), .Z(n30) );
  CLKBUF_X1 U51 ( .A(OP2[22]), .Z(n14) );
  CLKBUF_X1 U52 ( .A(OP2[26]), .Z(n15) );
  BUF_X2 U53 ( .A(OP2[1]), .Z(n16) );
  CLKBUF_X1 U54 ( .A(OP2[11]), .Z(n17) );
  BUF_X2 U55 ( .A(OP2[8]), .Z(n23) );
  CLKBUF_X1 U56 ( .A(OP2[10]), .Z(n19) );
  BUF_X2 U57 ( .A(OP2[2]), .Z(n38) );
  AND2_X1 U58 ( .A1(n55), .A2(n405), .ZN(n20) );
  NOR2_X1 U59 ( .A1(n20), .A2(n483), .ZN(n492) );
  INV_X2 U60 ( .A(n96), .ZN(n94) );
  AOI222_X1 U61 ( .A1(n47), .A2(n673), .B1(n657), .B2(n697), .C1(n238), .C2(
        n313), .ZN(n312) );
  AOI222_X1 U62 ( .A1(n375), .A2(n76), .B1(n373), .B2(n703), .C1(n689), .C2(
        n28), .ZN(n319) );
  AOI221_X1 U63 ( .B1(n364), .B2(n705), .C1(n153), .C2(n74), .A(n470), .ZN(
        n440) );
  AOI222_X1 U64 ( .A1(n47), .A2(n653), .B1(n663), .B2(n697), .C1(n238), .C2(
        n239), .ZN(n234) );
  AND2_X1 U65 ( .A1(n106), .A2(n107), .ZN(n21) );
  NAND2_X2 U66 ( .A1(n707), .A2(n704), .ZN(n460) );
  BUF_X2 U67 ( .A(OP2[5]), .Z(n22) );
  BUF_X2 U68 ( .A(OP2[14]), .Z(n24) );
  CLKBUF_X1 U69 ( .A(OP2[7]), .Z(n25) );
  INV_X2 U70 ( .A(n259), .ZN(n705) );
  CLKBUF_X1 U71 ( .A(OP2[9]), .Z(n27) );
  CLKBUF_X1 U72 ( .A(OP2[3]), .Z(n28) );
  AND2_X1 U73 ( .A1(n573), .A2(n62), .ZN(n29) );
  AND2_X1 U74 ( .A1(N189), .A2(n29), .ZN(n41) );
  INV_X1 U75 ( .A(n23), .ZN(n31) );
  INV_X1 U76 ( .A(n31), .ZN(n32) );
  CLKBUF_X1 U77 ( .A(OP2[20]), .Z(n33) );
  INV_X2 U78 ( .A(n58), .ZN(n91) );
  INV_X2 U79 ( .A(n96), .ZN(n93) );
  CLKBUF_X1 U80 ( .A(RES[30]), .Z(n34) );
  AOI211_X4 U81 ( .C1(n22), .C2(n57), .A(n212), .B(n215), .ZN(n130) );
  BUF_X1 U82 ( .A(n83), .Z(n35) );
  BUF_X1 U83 ( .A(n83), .Z(n36) );
  AND2_X2 U84 ( .A1(n709), .A2(n708), .ZN(n51) );
  CLKBUF_X1 U85 ( .A(n51), .Z(n83) );
  BUF_X1 U86 ( .A(n83), .Z(n88) );
  BUF_X1 U87 ( .A(n82), .Z(n86) );
  BUF_X1 U88 ( .A(n83), .Z(n87) );
  NAND2_X2 U89 ( .A1(n709), .A2(n708), .ZN(n337) );
  AOI222_X1 U90 ( .A1(n47), .A2(n671), .B1(n656), .B2(n697), .C1(n238), .C2(
        n299), .ZN(n298) );
  AOI221_X1 U91 ( .B1(n362), .B2(n705), .C1(n361), .C2(n74), .A(n672), .ZN(
        n305) );
  BUF_X2 U92 ( .A(n77), .Z(n79) );
  BUF_X1 U93 ( .A(n48), .Z(n77) );
  CLKBUF_X1 U94 ( .A(RES[31]), .Z(n37) );
  AOI222_X1 U95 ( .A1(n648), .A2(n47), .B1(n666), .B2(n697), .C1(n238), .C2(
        n581), .ZN(n579) );
  NAND2_X1 U96 ( .A1(n16), .A2(n63), .ZN(n240) );
  NAND2_X1 U97 ( .A1(n63), .A2(n50), .ZN(n257) );
  BUF_X2 U98 ( .A(OP2[0]), .Z(n63) );
  NAND2_X1 U99 ( .A1(N191), .A2(n7), .ZN(n106) );
  AND3_X1 U100 ( .A1(N189), .A2(n573), .A3(n62), .ZN(n39) );
  NAND3_X1 U101 ( .A1(n108), .A2(n105), .A3(n21), .ZN(RES[0]) );
  NOR2_X1 U102 ( .A1(n39), .A2(n4), .ZN(n40) );
  NOR2_X1 U103 ( .A1(n42), .A2(n41), .ZN(n108) );
  NAND2_X1 U104 ( .A1(n565), .A2(n9), .ZN(n42) );
  CLKBUF_X1 U105 ( .A(n105), .Z(n43) );
  CLKBUF_X1 U106 ( .A(n38), .Z(n44) );
  CLKBUF_X1 U107 ( .A(OP1[1]), .Z(n45) );
  INV_X1 U108 ( .A(n30), .ZN(n46) );
  INV_X2 U109 ( .A(n46), .ZN(n47) );
  AOI222_X4 U110 ( .A1(n47), .A2(n644), .B1(n664), .B2(n697), .C1(n238), .C2(
        n287), .ZN(n285) );
  AOI222_X4 U111 ( .A1(n47), .A2(n640), .B1(n665), .B2(n697), .C1(n238), .C2(
        n435), .ZN(n434) );
  AOI222_X4 U112 ( .A1(n47), .A2(n667), .B1(n255), .B2(n697), .C1(n238), .C2(
        n256), .ZN(n252) );
  AOI222_X4 U113 ( .A1(n47), .A2(n669), .B1(n655), .B2(n697), .C1(n238), .C2(
        n272), .ZN(n271) );
  AND2_X1 U114 ( .A1(n63), .A2(n50), .ZN(n48) );
  AND4_X1 U115 ( .A1(n40), .A2(n107), .A3(n106), .A4(n43), .ZN(n49) );
  INV_X1 U116 ( .A(OP2[1]), .ZN(n50) );
  NAND2_X1 U117 ( .A1(N193), .A2(n8), .ZN(n105) );
  BUF_X2 U118 ( .A(n48), .Z(n80) );
  BUF_X2 U119 ( .A(n48), .Z(n81) );
  CLKBUF_X1 U120 ( .A(n51), .Z(n82) );
  INV_X2 U121 ( .A(n97), .ZN(n92) );
  BUF_X1 U122 ( .A(n61), .Z(n68) );
  NAND2_X1 U123 ( .A1(N187), .A2(n68), .ZN(n52) );
  NAND2_X1 U124 ( .A1(N154), .A2(n66), .ZN(n53) );
  INV_X1 U125 ( .A(n502), .ZN(n54) );
  AND3_X1 U126 ( .A1(n53), .A2(n52), .A3(n54), .ZN(n503) );
  BUF_X1 U127 ( .A(n80), .Z(n78) );
  BUF_X1 U128 ( .A(n82), .Z(n84) );
  BUF_X1 U129 ( .A(n82), .Z(n85) );
  INV_X1 U130 ( .A(n395), .ZN(n615) );
  INV_X1 U131 ( .A(n460), .ZN(n703) );
  INV_X1 U132 ( .A(n219), .ZN(n699) );
  INV_X1 U133 ( .A(n236), .ZN(n698) );
  BUF_X1 U134 ( .A(n702), .Z(n75) );
  BUF_X1 U135 ( .A(n702), .Z(n74) );
  INV_X1 U136 ( .A(n97), .ZN(n95) );
  BUF_X1 U137 ( .A(n617), .Z(n71) );
  BUF_X1 U138 ( .A(n617), .Z(n72) );
  AND2_X1 U139 ( .A1(n73), .A2(n699), .ZN(n55) );
  BUF_X1 U140 ( .A(n702), .Z(n76) );
  BUF_X1 U141 ( .A(n617), .Z(n73) );
  NOR2_X1 U142 ( .A1(n147), .A2(n262), .ZN(n333) );
  NOR2_X1 U143 ( .A1(n262), .A2(n331), .ZN(n150) );
  NOR2_X1 U144 ( .A1(n147), .A2(n259), .ZN(n327) );
  NOR2_X1 U145 ( .A1(n259), .A2(n331), .ZN(n154) );
  NOR2_X1 U146 ( .A1(n147), .A2(n260), .ZN(n328) );
  NOR2_X1 U147 ( .A1(n331), .A2(n260), .ZN(n152) );
  INV_X1 U148 ( .A(n56), .ZN(n101) );
  INV_X1 U149 ( .A(n56), .ZN(n100) );
  INV_X1 U150 ( .A(n99), .ZN(n98) );
  INV_X1 U151 ( .A(n260), .ZN(n706) );
  NOR2_X1 U152 ( .A1(n389), .A2(n460), .ZN(n448) );
  NOR2_X1 U153 ( .A1(n526), .A2(n460), .ZN(n489) );
  NAND2_X1 U154 ( .A1(n6), .A2(n238), .ZN(n236) );
  NAND2_X1 U155 ( .A1(n238), .A2(n710), .ZN(n219) );
  INV_X1 U156 ( .A(n526), .ZN(n700) );
  INV_X1 U157 ( .A(OP2[0]), .ZN(n709) );
  INV_X1 U158 ( .A(n389), .ZN(n701) );
  NAND2_X1 U159 ( .A1(n124), .A2(n126), .ZN(n215) );
  BUF_X1 U160 ( .A(n59), .Z(n65) );
  BUF_X1 U161 ( .A(n59), .Z(n66) );
  INV_X1 U162 ( .A(n240), .ZN(n96) );
  INV_X1 U163 ( .A(n240), .ZN(n97) );
  BUF_X1 U164 ( .A(n59), .Z(n67) );
  INV_X1 U165 ( .A(n262), .ZN(n702) );
  INV_X1 U166 ( .A(n245), .ZN(n653) );
  INV_X1 U167 ( .A(n319), .ZN(n673) );
  INV_X1 U168 ( .A(n305), .ZN(n671) );
  INV_X1 U169 ( .A(n440), .ZN(n640) );
  INV_X1 U170 ( .A(n291), .ZN(n644) );
  INV_X1 U171 ( .A(n264), .ZN(n667) );
  INV_X1 U172 ( .A(n477), .ZN(n648) );
  NAND2_X1 U173 ( .A1(n127), .A2(n128), .ZN(n125) );
  OAI222_X1 U174 ( .A1(n257), .A2(n695), .B1(n89), .B2(n696), .C1(n337), .C2(
        n693), .ZN(n286) );
  OAI222_X1 U175 ( .A1(n257), .A2(n619), .B1(n89), .B2(n618), .C1(n337), .C2(
        n620), .ZN(n363) );
  OAI22_X1 U176 ( .A1(n337), .A2(n695), .B1(n257), .B2(n696), .ZN(n360) );
  AOI222_X1 U177 ( .A1(n237), .A2(n705), .B1(n387), .B2(n703), .C1(n391), .C2(
        n75), .ZN(n335) );
  AOI222_X1 U178 ( .A1(n360), .A2(n705), .B1(n361), .B2(n703), .C1(n362), .C2(
        n75), .ZN(n146) );
  AOI222_X1 U179 ( .A1(n286), .A2(n705), .B1(n402), .B2(n703), .C1(n404), .C2(
        n75), .ZN(n349) );
  AOI222_X1 U180 ( .A1(n375), .A2(n703), .B1(n705), .B2(n376), .C1(n377), .C2(
        n75), .ZN(n165) );
  OAI22_X1 U181 ( .A1(n337), .A2(n619), .B1(n257), .B2(n618), .ZN(n405) );
  AOI222_X1 U182 ( .A1(n392), .A2(n703), .B1(n705), .B2(n5), .C1(n393), .C2(
        n75), .ZN(n186) );
  AOI222_X1 U183 ( .A1(n392), .A2(n76), .B1(n183), .B2(n703), .C1(n654), .C2(
        n28), .ZN(n245) );
  INV_X1 U184 ( .A(n332), .ZN(n654) );
  AOI222_X1 U185 ( .A1(n378), .A2(n705), .B1(n169), .B2(n703), .C1(n379), .C2(
        n75), .ZN(n224) );
  AOI222_X1 U186 ( .A1(n363), .A2(n705), .B1(n153), .B2(n703), .C1(n364), .C2(
        n75), .ZN(n211) );
  AOI222_X1 U187 ( .A1(n405), .A2(n705), .B1(n406), .B2(n703), .C1(n407), .C2(
        n75), .ZN(n200) );
  INV_X1 U188 ( .A(n514), .ZN(n672) );
  AOI22_X1 U189 ( .A1(n703), .A2(n358), .B1(n706), .B2(n360), .ZN(n514) );
  OAI22_X1 U190 ( .A1(n460), .A2(n660), .B1(n260), .B2(n641), .ZN(n470) );
  INV_X1 U191 ( .A(n155), .ZN(n660) );
  OAI22_X1 U192 ( .A1(n460), .A2(n659), .B1(n260), .B2(n645), .ZN(n459) );
  INV_X1 U193 ( .A(n197), .ZN(n659) );
  AOI221_X1 U194 ( .B1(n404), .B2(n705), .C1(n402), .C2(n74), .A(n670), .ZN(
        n278) );
  INV_X1 U195 ( .A(n500), .ZN(n670) );
  AOI22_X1 U196 ( .A1(n703), .A2(n347), .B1(n706), .B2(n286), .ZN(n500) );
  AOI221_X1 U197 ( .B1(n391), .B2(n705), .C1(n387), .C2(n74), .A(n668), .ZN(
        n264) );
  INV_X1 U198 ( .A(n490), .ZN(n668) );
  AOI22_X1 U199 ( .A1(n703), .A2(n329), .B1(n706), .B2(n237), .ZN(n490) );
  AOI221_X1 U200 ( .B1(n379), .B2(n705), .C1(n169), .C2(n74), .A(n587), .ZN(
        n477) );
  OAI22_X1 U201 ( .A1(n460), .A2(n661), .B1(n649), .B2(n260), .ZN(n587) );
  INV_X1 U202 ( .A(n170), .ZN(n661) );
  INV_X1 U203 ( .A(n243), .ZN(n663) );
  AOI222_X1 U204 ( .A1(n182), .A2(n705), .B1(n184), .B2(n706), .C1(n185), .C2(
        n75), .ZN(n243) );
  INV_X1 U205 ( .A(n437), .ZN(n665) );
  AOI222_X1 U206 ( .A1(n156), .A2(n705), .B1(n151), .B2(n706), .C1(n210), .C2(
        n75), .ZN(n437) );
  INV_X1 U207 ( .A(n315), .ZN(n657) );
  AOI222_X1 U208 ( .A1(n316), .A2(n705), .B1(n317), .B2(n706), .C1(n318), .C2(
        n76), .ZN(n315) );
  INV_X1 U209 ( .A(n301), .ZN(n656) );
  AOI222_X1 U210 ( .A1(n302), .A2(n705), .B1(n303), .B2(n706), .C1(n304), .C2(
        n76), .ZN(n301) );
  AOI222_X1 U211 ( .A1(n275), .A2(n705), .B1(n276), .B2(n706), .C1(n277), .C2(
        n75), .ZN(n274) );
  AOI222_X1 U212 ( .A1(n171), .A2(n705), .B1(n168), .B2(n706), .C1(n683), .C2(
        n75), .ZN(n583) );
  INV_X1 U213 ( .A(n218), .ZN(n683) );
  OAI222_X1 U214 ( .A1(n658), .A2(n259), .B1(n662), .B2(n260), .C1(n261), .C2(
        n262), .ZN(n255) );
  INV_X1 U215 ( .A(n263), .ZN(n662) );
  NOR2_X1 U216 ( .A1(n696), .A2(n337), .ZN(n376) );
  OAI21_X1 U217 ( .B1(n22), .B2(n100), .A(n145), .ZN(n212) );
  OAI21_X1 U218 ( .B1(n2), .B2(n100), .A(n145), .ZN(n201) );
  OAI21_X1 U219 ( .B1(n25), .B2(n100), .A(n145), .ZN(n187) );
  OAI21_X1 U220 ( .B1(n32), .B2(n100), .A(n145), .ZN(n173) );
  OAI21_X1 U221 ( .B1(n27), .B2(n100), .A(n145), .ZN(n158) );
  AOI22_X1 U222 ( .A1(n237), .A2(n74), .B1(n391), .B2(n703), .ZN(n179) );
  AOI22_X1 U223 ( .A1(n360), .A2(n74), .B1(n362), .B2(n703), .ZN(n207) );
  AOI22_X1 U224 ( .A1(n286), .A2(n74), .B1(n404), .B2(n703), .ZN(n193) );
  NOR3_X1 U225 ( .A1(n147), .A2(n28), .A3(n223), .ZN(n222) );
  NOR3_X1 U226 ( .A1(n331), .A2(n28), .A3(n332), .ZN(n330) );
  AOI22_X1 U227 ( .A1(n363), .A2(n74), .B1(n364), .B2(n703), .ZN(n157) );
  AOI22_X1 U228 ( .A1(n405), .A2(n74), .B1(n407), .B2(n703), .ZN(n344) );
  AOI22_X1 U229 ( .A1(n378), .A2(n74), .B1(n379), .B2(n703), .ZN(n172) );
  NAND2_X1 U230 ( .A1(OP2[3]), .A2(n707), .ZN(n259) );
  OAI22_X1 U231 ( .A1(n234), .A2(n235), .B1(n691), .B2(n236), .ZN(n231) );
  INV_X1 U232 ( .A(n237), .ZN(n691) );
  OAI221_X1 U233 ( .B1(n95), .B2(n684), .C1(n90), .C2(n686), .A(n242), .ZN(
        n239) );
  OAI22_X1 U234 ( .A1(n434), .A2(n235), .B1(n694), .B2(n236), .ZN(n432) );
  INV_X1 U235 ( .A(n360), .ZN(n694) );
  OAI221_X1 U236 ( .B1(n95), .B2(n688), .C1(n90), .C2(n690), .A(n436), .ZN(
        n435) );
  OAI22_X1 U237 ( .A1(n285), .A2(n235), .B1(n692), .B2(n236), .ZN(n283) );
  INV_X1 U238 ( .A(n286), .ZN(n692) );
  OAI221_X1 U239 ( .B1(n95), .B2(n686), .C1(n89), .C2(n688), .A(n288), .ZN(
        n287) );
  OAI211_X1 U240 ( .C1(n193), .C2(n147), .A(n194), .B(n195), .ZN(n191) );
  AOI222_X1 U241 ( .A1(n150), .A2(n196), .B1(n152), .B2(n197), .C1(n154), .C2(
        n198), .ZN(n195) );
  AOI22_X1 U242 ( .A1(n700), .A2(n647), .B1(n699), .B2(n199), .ZN(n194) );
  INV_X1 U243 ( .A(n200), .ZN(n647) );
  OAI211_X1 U244 ( .C1(n179), .C2(n147), .A(n180), .B(n181), .ZN(n177) );
  AOI222_X1 U245 ( .A1(n150), .A2(n182), .B1(n152), .B2(n183), .C1(n154), .C2(
        n184), .ZN(n181) );
  AOI22_X1 U246 ( .A1(n700), .A2(n652), .B1(n699), .B2(n185), .ZN(n180) );
  INV_X1 U247 ( .A(n186), .ZN(n652) );
  NOR4_X1 U248 ( .A1(n599), .A2(OP2[23]), .A3(OP2[25]), .A4(OP2[24]), .ZN(n596) );
  NOR4_X1 U249 ( .A1(n601), .A2(n17), .A3(OP2[12]), .A4(OP2[10]), .ZN(n594) );
  NOR4_X1 U250 ( .A1(n600), .A2(OP2[16]), .A3(OP2[18]), .A4(OP2[17]), .ZN(n595) );
  AOI22_X1 U251 ( .A1(n150), .A2(n170), .B1(n699), .B2(n168), .ZN(n524) );
  AOI222_X1 U252 ( .A1(n154), .A2(n169), .B1(n489), .B2(n378), .C1(n152), .C2(
        n379), .ZN(n525) );
  AOI22_X1 U253 ( .A1(n150), .A2(n183), .B1(n699), .B2(n184), .ZN(n487) );
  AOI222_X1 U254 ( .A1(n154), .A2(n392), .B1(n489), .B2(n5), .C1(n152), .C2(
        n393), .ZN(n488) );
  AOI22_X1 U255 ( .A1(n150), .A2(n155), .B1(n699), .B2(n151), .ZN(n508) );
  AOI222_X1 U256 ( .A1(n154), .A2(n153), .B1(n489), .B2(n363), .C1(n152), .C2(
        n364), .ZN(n509) );
  AOI22_X1 U257 ( .A1(n150), .A2(n197), .B1(n699), .B2(n198), .ZN(n498) );
  AOI222_X1 U258 ( .A1(n154), .A2(n406), .B1(n489), .B2(n405), .C1(n152), .C2(
        n407), .ZN(n499) );
  AOI22_X1 U259 ( .A1(n333), .A2(n317), .B1(n698), .B2(n316), .ZN(n423) );
  AOI221_X1 U260 ( .B1(n327), .B2(n373), .C1(n328), .C2(n375), .A(n425), .ZN(
        n424) );
  NOR3_X1 U261 ( .A1(n389), .A2(n28), .A3(n223), .ZN(n425) );
  AOI22_X1 U262 ( .A1(n333), .A2(n329), .B1(n698), .B2(n263), .ZN(n446) );
  AOI222_X1 U263 ( .A1(n327), .A2(n387), .B1(n448), .B2(n237), .C1(n328), .C2(
        n391), .ZN(n447) );
  AOI222_X1 U264 ( .A1(n333), .A2(n275), .B1(n328), .B2(n347), .C1(n327), .C2(
        n276), .ZN(n346) );
  AOI22_X1 U265 ( .A1(n701), .A2(n677), .B1(n698), .B2(n277), .ZN(n345) );
  INV_X1 U266 ( .A(n349), .ZN(n677) );
  AOI22_X1 U267 ( .A1(n333), .A2(n358), .B1(n698), .B2(n303), .ZN(n467) );
  AOI222_X1 U268 ( .A1(n327), .A2(n361), .B1(n448), .B2(n360), .C1(n328), .C2(
        n362), .ZN(n468) );
  AOI22_X1 U269 ( .A1(n333), .A2(n373), .B1(n698), .B2(n317), .ZN(n478) );
  AOI222_X1 U270 ( .A1(n327), .A2(n375), .B1(n448), .B2(n376), .C1(n328), .C2(
        n377), .ZN(n479) );
  AOI22_X1 U271 ( .A1(n333), .A2(n347), .B1(n698), .B2(n276), .ZN(n456) );
  AOI222_X1 U272 ( .A1(n327), .A2(n402), .B1(n448), .B2(n286), .C1(n328), .C2(
        n404), .ZN(n457) );
  NAND2_X1 U273 ( .A1(n60), .A2(n580), .ZN(n235) );
  AOI22_X1 U274 ( .A1(n333), .A2(n334), .B1(n701), .B2(n675), .ZN(n325) );
  AOI221_X1 U275 ( .B1(n327), .B2(n263), .C1(n328), .C2(n329), .A(n330), .ZN(
        n326) );
  INV_X1 U276 ( .A(n335), .ZN(n675) );
  BUF_X1 U277 ( .A(n61), .Z(n69) );
  OAI211_X1 U278 ( .C1(n335), .C2(n147), .A(n536), .B(n537), .ZN(n534) );
  AOI22_X1 U279 ( .A1(n150), .A2(n184), .B1(n699), .B2(n182), .ZN(n536) );
  AOI221_X1 U280 ( .B1(n154), .B2(n183), .C1(n152), .C2(n392), .A(n538), .ZN(
        n537) );
  NOR3_X1 U281 ( .A1(n526), .A2(n28), .A3(n332), .ZN(n538) );
  OAI211_X1 U282 ( .C1(n207), .C2(n147), .A(n208), .B(n209), .ZN(n205) );
  AOI222_X1 U283 ( .A1(n150), .A2(n156), .B1(n152), .B2(n155), .C1(n154), .C2(
        n151), .ZN(n209) );
  AOI22_X1 U284 ( .A1(n700), .A2(n642), .B1(n699), .B2(n210), .ZN(n208) );
  INV_X1 U285 ( .A(n211), .ZN(n642) );
  AOI222_X1 U286 ( .A1(n333), .A2(n316), .B1(n328), .B2(n373), .C1(n327), .C2(
        n317), .ZN(n372) );
  AOI22_X1 U287 ( .A1(n701), .A2(n681), .B1(n698), .B2(n318), .ZN(n371) );
  INV_X1 U288 ( .A(n165), .ZN(n681) );
  OAI211_X1 U289 ( .C1(n218), .C2(n219), .A(n220), .B(n221), .ZN(n216) );
  AOI22_X1 U290 ( .A1(n150), .A2(n171), .B1(n700), .B2(n650), .ZN(n220) );
  AOI221_X1 U291 ( .B1(n154), .B2(n168), .C1(n152), .C2(n170), .A(n222), .ZN(
        n221) );
  INV_X1 U292 ( .A(n224), .ZN(n650) );
  OAI21_X1 U293 ( .B1(n17), .B2(n100), .A(n98), .ZN(n547) );
  OAI21_X1 U294 ( .B1(n100), .B2(OP2[10]), .A(n145), .ZN(n562) );
  OAI22_X1 U295 ( .A1(n389), .A2(n179), .B1(n236), .B2(n658), .ZN(n388) );
  AOI222_X1 U296 ( .A1(n333), .A2(n263), .B1(n328), .B2(n387), .C1(n327), .C2(
        n329), .ZN(n386) );
  OAI21_X1 U297 ( .B1(n28), .B2(n100), .A(n615), .ZN(n232) );
  OAI21_X1 U298 ( .B1(n16), .B2(n100), .A(n615), .ZN(n433) );
  BUF_X1 U299 ( .A(n61), .Z(n70) );
  OR4_X1 U300 ( .A1(OP2[19]), .A2(n33), .A3(OP2[21]), .A4(n14), .ZN(n600) );
  NOR4_X1 U301 ( .A1(n598), .A2(OP2[29]), .A3(n22), .A4(OP2[30]), .ZN(n597) );
  OR4_X1 U302 ( .A1(n2), .A2(n25), .A3(n23), .A4(n27), .ZN(n598) );
  INV_X1 U303 ( .A(OP2[3]), .ZN(n704) );
  AND2_X1 U304 ( .A1(n573), .A2(n574), .ZN(n56) );
  NAND2_X1 U305 ( .A1(n580), .A2(n573), .ZN(n126) );
  INV_X1 U306 ( .A(OP2[1]), .ZN(n708) );
  AND2_X1 U307 ( .A1(n60), .A2(n574), .ZN(n57) );
  AND2_X2 U308 ( .A1(n16), .A2(n709), .ZN(n58) );
  INV_X1 U309 ( .A(n334), .ZN(n658) );
  AND2_X1 U310 ( .A1(n62), .A2(n60), .ZN(n59) );
  INV_X1 U311 ( .A(n223), .ZN(n689) );
  AOI222_X1 U312 ( .A1(n333), .A2(n302), .B1(n328), .B2(n358), .C1(n327), .C2(
        n303), .ZN(n357) );
  AOI22_X1 U313 ( .A1(n701), .A2(n679), .B1(n698), .B2(n304), .ZN(n356) );
  INV_X1 U314 ( .A(n146), .ZN(n679) );
  NAND2_X1 U315 ( .A1(n593), .A2(n580), .ZN(n124) );
  AOI222_X1 U316 ( .A1(n333), .A2(n276), .B1(n328), .B2(n402), .C1(n327), .C2(
        n347), .ZN(n401) );
  AOI22_X1 U317 ( .A1(n701), .A2(n685), .B1(n698), .B2(n275), .ZN(n400) );
  INV_X1 U318 ( .A(n193), .ZN(n685) );
  OR3_X1 U319 ( .A1(n24), .A2(OP2[15]), .A3(n10), .ZN(n601) );
  OR3_X1 U320 ( .A1(OP2[27]), .A2(OP2[28]), .A3(n15), .ZN(n599) );
  OAI211_X1 U321 ( .C1(n146), .C2(n147), .A(n148), .B(n149), .ZN(n142) );
  AOI222_X1 U322 ( .A1(n150), .A2(n151), .B1(n152), .B2(n153), .C1(n154), .C2(
        n155), .ZN(n149) );
  AOI22_X1 U323 ( .A1(n700), .A2(n643), .B1(n699), .B2(n156), .ZN(n148) );
  INV_X1 U324 ( .A(n157), .ZN(n643) );
  AOI222_X1 U325 ( .A1(n333), .A2(n303), .B1(n328), .B2(n361), .C1(n327), .C2(
        n358), .ZN(n415) );
  AOI22_X1 U326 ( .A1(n701), .A2(n687), .B1(n698), .B2(n302), .ZN(n414) );
  INV_X1 U327 ( .A(n207), .ZN(n687) );
  OAI211_X1 U328 ( .C1(n165), .C2(n147), .A(n166), .B(n167), .ZN(n163) );
  AOI222_X1 U329 ( .A1(n150), .A2(n168), .B1(n152), .B2(n169), .C1(n154), .C2(
        n170), .ZN(n167) );
  AOI22_X1 U330 ( .A1(n700), .A2(n651), .B1(n699), .B2(n171), .ZN(n166) );
  INV_X1 U331 ( .A(n172), .ZN(n651) );
  OAI211_X1 U332 ( .C1(n349), .C2(n147), .A(n553), .B(n554), .ZN(n551) );
  AOI222_X1 U333 ( .A1(n150), .A2(n198), .B1(n152), .B2(n406), .C1(n154), .C2(
        n197), .ZN(n554) );
  AOI22_X1 U334 ( .A1(n700), .A2(n646), .B1(n699), .B2(n196), .ZN(n553) );
  INV_X1 U335 ( .A(n344), .ZN(n646) );
  INV_X1 U336 ( .A(n289), .ZN(n664) );
  AOI222_X1 U337 ( .A1(n196), .A2(n705), .B1(n198), .B2(n706), .C1(n199), .C2(
        n75), .ZN(n289) );
  OAI221_X1 U338 ( .B1(n95), .B2(n622), .C1(n89), .C2(n621), .A(n273), .ZN(
        n272) );
  INV_X1 U339 ( .A(n274), .ZN(n655) );
  INV_X1 U340 ( .A(n278), .ZN(n669) );
  AOI22_X1 U341 ( .A1(OP1[2]), .A2(n81), .B1(OP1[3]), .B2(n51), .ZN(n546) );
  INV_X1 U342 ( .A(n583), .ZN(n666) );
  AOI22_X1 U343 ( .A1(OP1[14]), .A2(n79), .B1(OP1[15]), .B2(n51), .ZN(n491) );
  AOI22_X1 U344 ( .A1(OP1[12]), .A2(n79), .B1(OP1[13]), .B2(n83), .ZN(n515) );
  AOI22_X1 U345 ( .A1(OP1[13]), .A2(n79), .B1(OP1[14]), .B2(n51), .ZN(n501) );
  AOI22_X1 U346 ( .A1(OP1[17]), .A2(n81), .B1(OP1[16]), .B2(n51), .ZN(n589) );
  AOI22_X1 U347 ( .A1(OP1[18]), .A2(n79), .B1(OP1[17]), .B2(n51), .ZN(n513) );
  OAI221_X1 U348 ( .B1(n625), .B2(n257), .C1(n626), .C2(n337), .A(n540), .ZN(
        n392) );
  AOI22_X1 U349 ( .A1(OP1[26]), .A2(n96), .B1(OP1[25]), .B2(n58), .ZN(n540) );
  OAI221_X1 U350 ( .B1(n93), .B2(n631), .C1(n90), .C2(n632), .A(n543), .ZN(
        n184) );
  AOI22_X1 U351 ( .A1(OP1[16]), .A2(n80), .B1(OP1[15]), .B2(n86), .ZN(n543) );
  OAI221_X1 U352 ( .B1(n94), .B2(n636), .C1(n90), .C2(n635), .A(n480), .ZN(
        n317) );
  AOI22_X1 U353 ( .A1(OP1[15]), .A2(n79), .B1(OP1[16]), .B2(n36), .ZN(n480) );
  OAI221_X1 U354 ( .B1(n93), .B2(n686), .C1(n90), .C2(n684), .A(n529), .ZN(
        n375) );
  AOI22_X1 U355 ( .A1(OP1[7]), .A2(n81), .B1(OP1[8]), .B2(n35), .ZN(n529) );
  OAI221_X1 U356 ( .B1(n93), .B2(n627), .C1(n90), .C2(n628), .A(n541), .ZN(
        n183) );
  AOI22_X1 U357 ( .A1(OP1[20]), .A2(n80), .B1(OP1[19]), .B2(n85), .ZN(n541) );
  AOI22_X1 U358 ( .A1(OP1[11]), .A2(n81), .B1(OP1[12]), .B2(n35), .ZN(n528) );
  AOI22_X1 U359 ( .A1(OP1[18]), .A2(n79), .B1(OP1[19]), .B2(n86), .ZN(n449) );
  OAI221_X1 U360 ( .B1(n94), .B2(n633), .C1(n90), .C2(n634), .A(n512), .ZN(
        n151) );
  AOI22_X1 U361 ( .A1(OP1[14]), .A2(n79), .B1(OP1[13]), .B2(n84), .ZN(n512) );
  AOI22_X1 U362 ( .A1(OP1[15]), .A2(n81), .B1(OP1[14]), .B2(n35), .ZN(n557) );
  AOI22_X1 U363 ( .A1(OP1[16]), .A2(n79), .B1(OP1[17]), .B2(n36), .ZN(n469) );
  OAI221_X1 U364 ( .B1(n94), .B2(n634), .C1(n90), .C2(n633), .A(n458), .ZN(
        n276) );
  AOI22_X1 U365 ( .A1(OP1[17]), .A2(n79), .B1(OP1[18]), .B2(n88), .ZN(n458) );
  AOI22_X1 U366 ( .A1(OP1[10]), .A2(n80), .B1(OP1[11]), .B2(n88), .ZN(n545) );
  OAI221_X1 U367 ( .B1(n93), .B2(n684), .C1(n90), .C2(n682), .A(n516), .ZN(
        n361) );
  AOI22_X1 U368 ( .A1(OP1[8]), .A2(n81), .B1(OP1[9]), .B2(n35), .ZN(n516) );
  OAI221_X1 U369 ( .B1(n94), .B2(n625), .C1(n89), .C2(n626), .A(n511), .ZN(
        n153) );
  AOI22_X1 U370 ( .A1(OP1[22]), .A2(n79), .B1(OP1[21]), .B2(n87), .ZN(n511) );
  OAI221_X1 U371 ( .B1(n94), .B2(n624), .C1(n625), .C2(n89), .A(n556), .ZN(
        n406) );
  AOI22_X1 U372 ( .A1(n80), .A2(OP1[23]), .B1(n36), .B2(OP1[22]), .ZN(n556) );
  AOI22_X1 U373 ( .A1(OP1[9]), .A2(n80), .B1(OP1[10]), .B2(n84), .ZN(n561) );
  AOI22_X1 U374 ( .A1(OP1[6]), .A2(n81), .B1(OP1[7]), .B2(n87), .ZN(n544) );
  AOI22_X1 U375 ( .A1(OP1[26]), .A2(n79), .B1(OP1[25]), .B2(n87), .ZN(n510) );
  OAI221_X1 U376 ( .B1(n93), .B2(n693), .C1(n90), .C2(n690), .A(n517), .ZN(
        n362) );
  AOI22_X1 U377 ( .A1(OP1[4]), .A2(n80), .B1(OP1[5]), .B2(n87), .ZN(n517) );
  AOI22_X1 U378 ( .A1(OP1[27]), .A2(n81), .B1(OP1[26]), .B2(n86), .ZN(n559) );
  AOI22_X1 U379 ( .A1(OP1[5]), .A2(n80), .B1(OP1[6]), .B2(n87), .ZN(n560) );
  OAI221_X1 U380 ( .B1(n257), .B2(n628), .C1(n627), .C2(n337), .A(n403), .ZN(
        n275) );
  AOI22_X1 U381 ( .A1(OP1[19]), .A2(n96), .B1(OP1[20]), .B2(n58), .ZN(n403) );
  OAI221_X1 U382 ( .B1(n95), .B2(n631), .C1(n89), .C2(n630), .A(n416), .ZN(
        n302) );
  AOI22_X1 U383 ( .A1(OP1[20]), .A2(n78), .B1(OP1[21]), .B2(n35), .ZN(n416) );
  AOI22_X1 U384 ( .A1(OP1[19]), .A2(n78), .B1(OP1[20]), .B2(n85), .ZN(n426) );
  OAI221_X1 U385 ( .B1(n93), .B2(n635), .C1(n90), .C2(n636), .A(n542), .ZN(
        n182) );
  AOI22_X1 U386 ( .A1(OP1[12]), .A2(n81), .B1(OP1[11]), .B2(n88), .ZN(n542) );
  AOI22_X1 U387 ( .A1(OP1[10]), .A2(n79), .B1(OP1[9]), .B2(n86), .ZN(n439) );
  AOI22_X1 U388 ( .A1(OP1[11]), .A2(n80), .B1(OP1[10]), .B2(n87), .ZN(n558) );
  OAI221_X1 U389 ( .B1(n93), .B2(n619), .C1(n90), .C2(n620), .A(n539), .ZN(
        n393) );
  AOI22_X1 U390 ( .A1(OP1[28]), .A2(n81), .B1(OP1[27]), .B2(n51), .ZN(n539) );
  OAI221_X1 U391 ( .B1(n257), .B2(n627), .C1(n626), .C2(n337), .A(n390), .ZN(
        n334) );
  AOI22_X1 U392 ( .A1(OP1[20]), .A2(n96), .B1(OP1[21]), .B2(n58), .ZN(n390) );
  OAI221_X1 U393 ( .B1(n626), .B2(n257), .C1(n625), .C2(n337), .A(n374), .ZN(
        n318) );
  AOI22_X1 U394 ( .A1(OP1[21]), .A2(n97), .B1(OP1[22]), .B2(n58), .ZN(n374) );
  OAI221_X1 U395 ( .B1(n625), .B2(n257), .C1(n337), .C2(n624), .A(n359), .ZN(
        n304) );
  AOI22_X1 U396 ( .A1(OP1[22]), .A2(n97), .B1(OP1[23]), .B2(n58), .ZN(n359) );
  OAI221_X1 U397 ( .B1(n95), .B2(n626), .C1(n625), .C2(n89), .A(n348), .ZN(
        n277) );
  AOI22_X1 U398 ( .A1(OP1[25]), .A2(n78), .B1(OP1[26]), .B2(n36), .ZN(n348) );
  OAI221_X1 U399 ( .B1(n95), .B2(n676), .C1(n89), .C2(n678), .A(n244), .ZN(
        n185) );
  AOI22_X1 U400 ( .A1(OP1[8]), .A2(n78), .B1(OP1[7]), .B2(n85), .ZN(n244) );
  OAI221_X1 U401 ( .B1(n95), .B2(n680), .C1(n89), .C2(n682), .A(n438), .ZN(
        n210) );
  AOI22_X1 U402 ( .A1(OP1[6]), .A2(n78), .B1(OP1[5]), .B2(n36), .ZN(n438) );
  OAI221_X1 U403 ( .B1(n95), .B2(n678), .C1(n89), .C2(n680), .A(n290), .ZN(
        n199) );
  AOI22_X1 U404 ( .A1(OP1[7]), .A2(n78), .B1(OP1[6]), .B2(n84), .ZN(n290) );
  NOR2_X1 U405 ( .A1(n711), .A2(ALU_OP[2]), .ZN(n580) );
  AOI21_X1 U406 ( .B1(OP1[28]), .B2(n97), .A(n5), .ZN(n258) );
  AOI221_X1 U407 ( .B1(n96), .B2(OP1[24]), .C1(n58), .C2(OP1[25]), .A(n336), 
        .ZN(n261) );
  OAI22_X1 U408 ( .A1(n623), .A2(n257), .B1(n622), .B2(n337), .ZN(n336) );
  AOI221_X1 U409 ( .B1(n97), .B2(OP1[7]), .C1(n58), .C2(OP1[6]), .A(n584), 
        .ZN(n218) );
  OAI22_X1 U410 ( .A1(n686), .A2(n257), .B1(n688), .B2(n337), .ZN(n584) );
  OAI221_X1 U411 ( .B1(n95), .B2(n624), .C1(n89), .C2(n623), .A(n314), .ZN(
        n313) );
  AOI22_X1 U412 ( .A1(OP1[27]), .A2(n78), .B1(OP1[28]), .B2(n84), .ZN(n314) );
  OAI221_X1 U413 ( .B1(n95), .B2(n623), .C1(n89), .C2(n622), .A(n300), .ZN(
        n299) );
  AOI22_X1 U414 ( .A1(OP1[28]), .A2(n78), .B1(OP1[29]), .B2(n51), .ZN(n300) );
  OAI221_X1 U415 ( .B1(n94), .B2(n626), .C1(n89), .C2(n627), .A(n590), .ZN(
        n169) );
  AOI22_X1 U416 ( .A1(OP1[21]), .A2(n78), .B1(OP1[20]), .B2(n82), .ZN(n590) );
  AOI22_X1 U417 ( .A1(OP1[4]), .A2(n81), .B1(OP1[3]), .B2(n35), .ZN(n242) );
  OAI221_X1 U418 ( .B1(n257), .B2(n624), .C1(n625), .C2(n337), .A(n591), .ZN(
        n379) );
  AOI22_X1 U419 ( .A1(OP1[27]), .A2(n96), .B1(OP1[26]), .B2(n58), .ZN(n591) );
  AOI22_X1 U420 ( .A1(OP1[9]), .A2(n80), .B1(OP1[8]), .B2(n51), .ZN(n586) );
  OAI221_X1 U421 ( .B1(n93), .B2(n695), .C1(n90), .C2(n693), .A(n527), .ZN(
        n377) );
  AOI22_X1 U422 ( .A1(OP1[3]), .A2(n81), .B1(OP1[4]), .B2(n51), .ZN(n527) );
  AOI22_X1 U423 ( .A1(OP1[3]), .A2(n78), .B1(OP1[2]), .B2(n36), .ZN(n288) );
  AOI22_X1 U424 ( .A1(OP1[29]), .A2(n77), .B1(OP1[28]), .B2(n51), .ZN(n588) );
  AOI22_X1 U425 ( .A1(OP1[19]), .A2(n80), .B1(OP1[18]), .B2(n51), .ZN(n555) );
  AOI22_X1 U426 ( .A1(OP1[13]), .A2(n80), .B1(OP1[12]), .B2(n83), .ZN(n585) );
  INV_X1 U427 ( .A(OP1[5]), .ZN(n686) );
  INV_X1 U428 ( .A(OP1[4]), .ZN(n688) );
  INV_X1 U429 ( .A(n45), .ZN(n695) );
  INV_X1 U430 ( .A(OP1[11]), .ZN(n674) );
  INV_X1 U431 ( .A(OP1[10]), .ZN(n676) );
  INV_X1 U433 ( .A(OP1[8]), .ZN(n680) );
  INV_X1 U434 ( .A(OP1[9]), .ZN(n678) );
  INV_X1 U435 ( .A(OP1[7]), .ZN(n682) );
  INV_X1 U436 ( .A(OP1[6]), .ZN(n684) );
  INV_X1 U437 ( .A(OP1[3]), .ZN(n690) );
  NOR2_X1 U438 ( .A1(n638), .A2(ALU_OP[0]), .ZN(n573) );
  AOI22_X1 U439 ( .A1(OP1[2]), .A2(n78), .B1(n45), .B2(n85), .ZN(n436) );
  AOI22_X1 U440 ( .A1(OP1[29]), .A2(n78), .B1(OP1[30]), .B2(n86), .ZN(n273) );
  AOI21_X1 U441 ( .B1(OP1[3]), .B2(n97), .A(n376), .ZN(n582) );
  INV_X1 U443 ( .A(OP1[2]), .ZN(n693) );
  OAI21_X1 U444 ( .B1(OP1[4]), .B2(n100), .A(n98), .ZN(n217) );
  OAI21_X1 U445 ( .B1(OP1[5]), .B2(n100), .A(n145), .ZN(n206) );
  OAI21_X1 U446 ( .B1(OP1[6]), .B2(n101), .A(n145), .ZN(n192) );
  OAI21_X1 U447 ( .B1(OP1[7]), .B2(n100), .A(n145), .ZN(n178) );
  OAI21_X1 U448 ( .B1(OP1[8]), .B2(n100), .A(n145), .ZN(n164) );
  OAI21_X1 U449 ( .B1(OP1[9]), .B2(n100), .A(n145), .ZN(n143) );
  OAI21_X1 U450 ( .B1(OP1[10]), .B2(n100), .A(n98), .ZN(n552) );
  INV_X1 U451 ( .A(n18), .ZN(n696) );
  OAI21_X1 U452 ( .B1(OP1[11]), .B2(n100), .A(n145), .ZN(n535) );
  AND2_X1 U453 ( .A1(n102), .A2(n638), .ZN(n60) );
  AND2_X1 U454 ( .A1(ALU_OP[2]), .A2(n711), .ZN(n574) );
  AND3_X1 U455 ( .A1(ALU_OP[0]), .A2(n638), .A3(n62), .ZN(n61) );
  AND2_X1 U456 ( .A1(ALU_OP[0]), .A2(ALU_OP[1]), .ZN(n593) );
  AOI21_X1 U457 ( .B1(n18), .B2(n576), .A(n577), .ZN(n565) );
  OAI211_X1 U458 ( .C1(n63), .C2(n100), .A(n592), .B(n616), .ZN(n576) );
  INV_X1 U459 ( .A(ALU_OP[3]), .ZN(n711) );
  NOR2_X1 U460 ( .A1(ALU_OP[2]), .A2(ALU_OP[3]), .ZN(n62) );
  OAI22_X1 U461 ( .A1(n639), .A2(n124), .B1(n125), .B2(n126), .ZN(ZERO) );
  INV_X1 U462 ( .A(n125), .ZN(n639) );
  OAI21_X1 U463 ( .B1(n44), .B2(n100), .A(n615), .ZN(n284) );
  AOI22_X1 U464 ( .A1(n377), .A2(n707), .B1(n44), .B2(n376), .ZN(n223) );
  AOI22_X1 U465 ( .A1(n707), .A2(n393), .B1(n44), .B2(n5), .ZN(n332) );
  NAND2_X1 U466 ( .A1(n38), .A2(OP2[3]), .ZN(n260) );
  NAND2_X1 U467 ( .A1(n38), .A2(n704), .ZN(n262) );
  INV_X1 U468 ( .A(n38), .ZN(n707) );
  OAI21_X1 U469 ( .B1(n47), .B2(n100), .A(n98), .ZN(n225) );
  NAND2_X1 U470 ( .A1(n47), .A2(n710), .ZN(n526) );
  NAND2_X1 U471 ( .A1(n6), .A2(n47), .ZN(n389) );
  NOR2_X1 U472 ( .A1(n460), .A2(n47), .ZN(n238) );
  INV_X1 U473 ( .A(n30), .ZN(n697) );
  INV_X1 U474 ( .A(n57), .ZN(n64) );
  INV_X1 U475 ( .A(n145), .ZN(n99) );
  INV_X1 U476 ( .A(ALU_OP[1]), .ZN(n638) );
  NAND3_X1 U477 ( .A1(n574), .A2(ALU_OP[0]), .A3(n638), .ZN(n145) );
  NAND2_X1 U478 ( .A1(n709), .A2(n696), .ZN(n104) );
  INV_X1 U479 ( .A(ALU_OP[0]), .ZN(n102) );
  NOR3_X1 U480 ( .A1(n709), .A2(n64), .A3(n696), .ZN(n103) );
  AOI221_X1 U481 ( .B1(n104), .B2(n99), .C1(N123), .C2(n65), .A(n103), .ZN(
        n107) );
  NAND4_X1 U482 ( .A1(n596), .A2(n597), .A3(n594), .A4(n595), .ZN(n578) );
  MUX2_X1 U483 ( .A(n64), .B(n101), .S(n695), .Z(n109) );
  AOI21_X1 U484 ( .B1(n109), .B2(n98), .A(n708), .ZN(n110) );
  AOI221_X1 U485 ( .B1(N157), .B2(n68), .C1(N124), .C2(n65), .A(n110), .ZN(
        n112) );
  INV_X1 U486 ( .A(n578), .ZN(n617) );
  AOI22_X1 U487 ( .A1(n432), .A2(n72), .B1(n45), .B2(n433), .ZN(n111) );
  NAND2_X1 U488 ( .A1(n111), .A2(n112), .ZN(RES[1]) );
  MUX2_X1 U489 ( .A(n64), .B(n101), .S(n693), .Z(n113) );
  AOI21_X1 U490 ( .B1(n113), .B2(n98), .A(n707), .ZN(n114) );
  AOI221_X1 U491 ( .B1(N158), .B2(n69), .C1(N125), .C2(n65), .A(n114), .ZN(
        n116) );
  AOI22_X1 U492 ( .A1(n283), .A2(n72), .B1(OP1[2]), .B2(n284), .ZN(n115) );
  NAND2_X1 U493 ( .A1(n116), .A2(n115), .ZN(RES[2]) );
  MUX2_X1 U494 ( .A(n64), .B(n101), .S(n690), .Z(n117) );
  AOI21_X1 U495 ( .B1(n117), .B2(n98), .A(n704), .ZN(n118) );
  AOI221_X1 U496 ( .B1(N159), .B2(n69), .C1(N126), .C2(n65), .A(n118), .ZN(
        n120) );
  AOI22_X1 U497 ( .A1(n231), .A2(n73), .B1(OP1[3]), .B2(n232), .ZN(n119) );
  NAND2_X1 U498 ( .A1(n120), .A2(n119), .ZN(RES[3]) );
  NOR2_X1 U499 ( .A1(n688), .A2(n121), .ZN(n122) );
  AOI221_X1 U500 ( .B1(N160), .B2(n69), .C1(N127), .C2(n65), .A(n122), .ZN(
        n129) );
  AOI22_X1 U501 ( .A1(n216), .A2(n73), .B1(n217), .B2(n47), .ZN(n123) );
  NAND2_X1 U502 ( .A1(n129), .A2(n123), .ZN(RES[4]) );
  NOR2_X1 U503 ( .A1(n686), .A2(n130), .ZN(n131) );
  AOI221_X1 U504 ( .B1(N161), .B2(n69), .C1(N128), .C2(n65), .A(n131), .ZN(
        n133) );
  AOI22_X1 U505 ( .A1(n205), .A2(n72), .B1(n206), .B2(n22), .ZN(n132) );
  NAND2_X1 U506 ( .A1(n133), .A2(n132), .ZN(RES[5]) );
  NOR2_X1 U507 ( .A1(n684), .A2(n134), .ZN(n135) );
  AOI221_X1 U508 ( .B1(N162), .B2(n69), .C1(N129), .C2(n65), .A(n135), .ZN(
        n137) );
  AOI22_X1 U509 ( .A1(n191), .A2(n72), .B1(n192), .B2(n2), .ZN(n136) );
  NAND2_X1 U510 ( .A1(n137), .A2(n136), .ZN(RES[6]) );
  AOI211_X1 U511 ( .C1(n25), .C2(n57), .A(n187), .B(n215), .ZN(n138) );
  NOR2_X1 U512 ( .A1(n682), .A2(n138), .ZN(n139) );
  AOI221_X1 U513 ( .B1(N163), .B2(n68), .C1(N130), .C2(n65), .A(n139), .ZN(
        n141) );
  AOI22_X1 U514 ( .A1(n177), .A2(n72), .B1(n178), .B2(n25), .ZN(n140) );
  NAND2_X1 U515 ( .A1(n141), .A2(n140), .ZN(RES[7]) );
  NOR2_X1 U516 ( .A1(n680), .A2(n144), .ZN(n159) );
  AOI221_X1 U517 ( .B1(N164), .B2(n68), .C1(N131), .C2(n65), .A(n159), .ZN(
        n161) );
  AOI22_X1 U518 ( .A1(n163), .A2(n72), .B1(n164), .B2(n32), .ZN(n160) );
  NAND2_X1 U519 ( .A1(n161), .A2(n160), .ZN(RES[8]) );
  AOI211_X1 U520 ( .C1(n27), .C2(n57), .A(n158), .B(n215), .ZN(n162) );
  NOR2_X1 U521 ( .A1(n678), .A2(n162), .ZN(n174) );
  AOI221_X1 U522 ( .B1(N165), .B2(n68), .C1(N132), .C2(n65), .A(n174), .ZN(
        n176) );
  AOI22_X1 U523 ( .A1(n142), .A2(n72), .B1(n143), .B2(n27), .ZN(n175) );
  NAND2_X1 U524 ( .A1(n176), .A2(n175), .ZN(RES[9]) );
  NOR2_X1 U525 ( .A1(n676), .A2(n188), .ZN(n189) );
  AOI221_X1 U526 ( .B1(N166), .B2(n68), .C1(N133), .C2(n65), .A(n189), .ZN(
        n202) );
  AOI22_X1 U527 ( .A1(n551), .A2(n72), .B1(n552), .B2(n19), .ZN(n190) );
  NAND2_X1 U528 ( .A1(n202), .A2(n190), .ZN(RES[10]) );
  AOI211_X1 U529 ( .C1(n17), .C2(n57), .A(n547), .B(n215), .ZN(n203) );
  NOR2_X1 U530 ( .A1(n674), .A2(n203), .ZN(n204) );
  AOI221_X1 U531 ( .B1(N167), .B2(n68), .C1(N134), .C2(n65), .A(n204), .ZN(
        n214) );
  AOI22_X1 U532 ( .A1(n534), .A2(n72), .B1(n535), .B2(n17), .ZN(n213) );
  NAND2_X1 U533 ( .A1(n214), .A2(n213), .ZN(RES[11]) );
  OAI21_X1 U534 ( .B1(OP1[12]), .B2(n100), .A(n98), .ZN(n229) );
  OAI211_X1 U535 ( .C1(n319), .C2(n147), .A(n524), .B(n525), .ZN(n228) );
  INV_X1 U536 ( .A(n215), .ZN(n616) );
  NAND2_X1 U537 ( .A1(n616), .A2(n145), .ZN(n395) );
  MUX2_X1 U538 ( .A(n101), .B(n64), .S(OP2[12]), .Z(n226) );
  INV_X1 U539 ( .A(OP1[12]), .ZN(n637) );
  AOI21_X1 U540 ( .B1(n615), .B2(n226), .A(n637), .ZN(n227) );
  AOI221_X1 U541 ( .B1(OP2[12]), .B2(n229), .C1(n228), .C2(n72), .A(n227), 
        .ZN(n233) );
  AOI22_X1 U542 ( .A1(N135), .A2(n66), .B1(N168), .B2(n69), .ZN(n230) );
  NAND2_X1 U543 ( .A1(n233), .A2(n230), .ZN(RES[12]) );
  OAI21_X1 U544 ( .B1(OP1[13]), .B2(n101), .A(n145), .ZN(n248) );
  OAI211_X1 U545 ( .C1(n305), .C2(n147), .A(n508), .B(n509), .ZN(n247) );
  MUX2_X1 U546 ( .A(n101), .B(n64), .S(n10), .Z(n241) );
  INV_X1 U547 ( .A(OP1[13]), .ZN(n636) );
  AOI21_X1 U548 ( .B1(n615), .B2(n241), .A(n636), .ZN(n246) );
  AOI221_X1 U549 ( .B1(n10), .B2(n248), .C1(n247), .C2(n72), .A(n246), .ZN(
        n250) );
  AOI22_X1 U550 ( .A1(N136), .A2(n67), .B1(N169), .B2(n69), .ZN(n249) );
  NAND2_X1 U551 ( .A1(n250), .A2(n249), .ZN(RES[13]) );
  OAI21_X1 U552 ( .B1(OP1[14]), .B2(n100), .A(n145), .ZN(n265) );
  OAI211_X1 U553 ( .C1(n278), .C2(n147), .A(n498), .B(n499), .ZN(n254) );
  MUX2_X1 U554 ( .A(n101), .B(n64), .S(n24), .Z(n251) );
  INV_X1 U555 ( .A(OP1[14]), .ZN(n635) );
  AOI21_X1 U556 ( .B1(n615), .B2(n251), .A(n635), .ZN(n253) );
  AOI221_X1 U557 ( .B1(n24), .B2(n265), .C1(n254), .C2(n71), .A(n253), .ZN(
        n267) );
  AOI22_X1 U558 ( .A1(N137), .A2(n67), .B1(N170), .B2(n69), .ZN(n266) );
  NAND2_X1 U559 ( .A1(n267), .A2(n266), .ZN(RES[14]) );
  OAI21_X1 U560 ( .B1(OP1[15]), .B2(n100), .A(n145), .ZN(n279) );
  OAI211_X1 U561 ( .C1(n264), .C2(n147), .A(n487), .B(n488), .ZN(n270) );
  MUX2_X1 U562 ( .A(n101), .B(n64), .S(OP2[15]), .Z(n268) );
  INV_X1 U563 ( .A(OP1[15]), .ZN(n634) );
  AOI21_X1 U564 ( .B1(n615), .B2(n268), .A(n634), .ZN(n269) );
  AOI221_X1 U565 ( .B1(OP2[15]), .B2(n279), .C1(n270), .C2(n72), .A(n269), 
        .ZN(n281) );
  AOI22_X1 U566 ( .A1(N138), .A2(n67), .B1(N171), .B2(n69), .ZN(n280) );
  NAND2_X1 U567 ( .A1(n281), .A2(n280), .ZN(RES[15]) );
  OAI21_X1 U568 ( .B1(OP1[16]), .B2(n100), .A(n98), .ZN(n294) );
  OAI211_X1 U569 ( .C1(n26), .C2(n331), .A(n478), .B(n479), .ZN(n293) );
  MUX2_X1 U570 ( .A(n101), .B(n64), .S(OP2[16]), .Z(n282) );
  INV_X1 U571 ( .A(OP1[16]), .ZN(n633) );
  AOI21_X1 U572 ( .B1(n615), .B2(n282), .A(n633), .ZN(n292) );
  AOI221_X1 U573 ( .B1(OP2[16]), .B2(n294), .C1(n293), .C2(n71), .A(n292), 
        .ZN(n296) );
  AOI22_X1 U574 ( .A1(N139), .A2(n67), .B1(N172), .B2(n69), .ZN(n295) );
  NAND2_X1 U575 ( .A1(n296), .A2(n295), .ZN(RES[16]) );
  OAI21_X1 U576 ( .B1(OP1[17]), .B2(n100), .A(n145), .ZN(n308) );
  OAI211_X1 U577 ( .C1(n440), .C2(n331), .A(n467), .B(n468), .ZN(n307) );
  MUX2_X1 U578 ( .A(n101), .B(n64), .S(OP2[17]), .Z(n297) );
  INV_X1 U579 ( .A(OP1[17]), .ZN(n632) );
  AOI21_X1 U580 ( .B1(n615), .B2(n297), .A(n632), .ZN(n306) );
  AOI221_X1 U581 ( .B1(OP2[17]), .B2(n308), .C1(n307), .C2(n71), .A(n306), 
        .ZN(n310) );
  AOI22_X1 U582 ( .A1(N140), .A2(n66), .B1(N173), .B2(n69), .ZN(n309) );
  NAND2_X1 U583 ( .A1(n310), .A2(n309), .ZN(RES[17]) );
  OAI21_X1 U584 ( .B1(OP1[18]), .B2(n100), .A(n145), .ZN(n322) );
  OAI211_X1 U585 ( .C1(n291), .C2(n331), .A(n456), .B(n457), .ZN(n321) );
  MUX2_X1 U586 ( .A(n101), .B(n64), .S(OP2[18]), .Z(n311) );
  INV_X1 U587 ( .A(OP1[18]), .ZN(n631) );
  AOI21_X1 U588 ( .B1(n615), .B2(n311), .A(n631), .ZN(n320) );
  AOI221_X1 U589 ( .B1(OP2[18]), .B2(n322), .C1(n321), .C2(n71), .A(n320), 
        .ZN(n324) );
  AOI22_X1 U590 ( .A1(N141), .A2(n67), .B1(N174), .B2(n69), .ZN(n323) );
  NAND2_X1 U591 ( .A1(n324), .A2(n323), .ZN(RES[18]) );
  OAI21_X1 U592 ( .B1(OP1[19]), .B2(n101), .A(n145), .ZN(n341) );
  OAI211_X1 U593 ( .C1(n245), .C2(n331), .A(n446), .B(n447), .ZN(n340) );
  MUX2_X1 U594 ( .A(n101), .B(n64), .S(OP2[19]), .Z(n338) );
  INV_X1 U595 ( .A(OP1[19]), .ZN(n630) );
  AOI21_X1 U596 ( .B1(n615), .B2(n338), .A(n630), .ZN(n339) );
  AOI221_X1 U597 ( .B1(OP2[19]), .B2(n341), .C1(n340), .C2(n71), .A(n339), 
        .ZN(n343) );
  AOI22_X1 U598 ( .A1(N142), .A2(n67), .B1(N175), .B2(n70), .ZN(n342) );
  NAND2_X1 U599 ( .A1(n343), .A2(n342), .ZN(RES[19]) );
  OAI21_X1 U600 ( .B1(OP1[20]), .B2(n101), .A(n98), .ZN(n353) );
  OAI211_X1 U601 ( .C1(n224), .C2(n331), .A(n423), .B(n424), .ZN(n352) );
  MUX2_X1 U602 ( .A(n101), .B(n64), .S(n33), .Z(n350) );
  INV_X1 U603 ( .A(OP1[20]), .ZN(n629) );
  AOI21_X1 U604 ( .B1(n615), .B2(n350), .A(n629), .ZN(n351) );
  AOI221_X1 U605 ( .B1(n33), .B2(n353), .C1(n352), .C2(n71), .A(n351), .ZN(
        n355) );
  AOI22_X1 U606 ( .A1(N143), .A2(n67), .B1(N176), .B2(n70), .ZN(n354) );
  NAND2_X1 U607 ( .A1(n355), .A2(n354), .ZN(RES[20]) );
  OAI21_X1 U608 ( .B1(OP1[21]), .B2(n101), .A(n98), .ZN(n368) );
  OAI211_X1 U609 ( .C1(n211), .C2(n331), .A(n414), .B(n415), .ZN(n367) );
  MUX2_X1 U610 ( .A(n101), .B(n64), .S(OP2[21]), .Z(n365) );
  INV_X1 U611 ( .A(OP1[21]), .ZN(n628) );
  AOI21_X1 U612 ( .B1(n615), .B2(n365), .A(n628), .ZN(n366) );
  AOI221_X1 U613 ( .B1(OP2[21]), .B2(n368), .C1(n367), .C2(n71), .A(n366), 
        .ZN(n370) );
  AOI22_X1 U614 ( .A1(N144), .A2(n66), .B1(N177), .B2(n70), .ZN(n369) );
  NAND2_X1 U615 ( .A1(n370), .A2(n369), .ZN(RES[21]) );
  OAI21_X1 U616 ( .B1(OP1[22]), .B2(n101), .A(n98), .ZN(n383) );
  OAI211_X1 U617 ( .C1(n200), .C2(n331), .A(n400), .B(n401), .ZN(n382) );
  MUX2_X1 U618 ( .A(n101), .B(n64), .S(n14), .Z(n380) );
  INV_X1 U619 ( .A(OP1[22]), .ZN(n627) );
  AOI21_X1 U620 ( .B1(n615), .B2(n380), .A(n627), .ZN(n381) );
  AOI221_X1 U621 ( .B1(n14), .B2(n383), .C1(n382), .C2(n71), .A(n381), .ZN(
        n385) );
  AOI22_X1 U622 ( .A1(N145), .A2(n66), .B1(N178), .B2(n70), .ZN(n384) );
  NAND2_X1 U623 ( .A1(n385), .A2(n384), .ZN(RES[22]) );
  INV_X1 U624 ( .A(OP1[23]), .ZN(n626) );
  AOI21_X1 U625 ( .B1(n56), .B2(n626), .A(n99), .ZN(n408) );
  INV_X1 U628 ( .A(OP2[23]), .ZN(n399) );
  OAI21_X1 U629 ( .B1(n186), .B2(n331), .A(n386), .ZN(n394) );
  OAI21_X1 U630 ( .B1(n388), .B2(n394), .A(n73), .ZN(n398) );
  MUX2_X1 U631 ( .A(n56), .B(n57), .S(OP2[23]), .Z(n396) );
  OAI21_X1 U632 ( .B1(n396), .B2(n395), .A(OP1[23]), .ZN(n397) );
  OAI211_X1 U633 ( .C1(n408), .C2(n399), .A(n398), .B(n397), .ZN(n409) );
  AOI221_X1 U634 ( .B1(N146), .B2(n67), .C1(N179), .C2(n68), .A(n409), .ZN(
        n548) );
  INV_X1 U635 ( .A(n548), .ZN(RES[23]) );
  OAI21_X1 U636 ( .B1(OP1[24]), .B2(n101), .A(n98), .ZN(n413) );
  OAI211_X1 U637 ( .C1(n172), .C2(n331), .A(n371), .B(n372), .ZN(n412) );
  MUX2_X1 U638 ( .A(n101), .B(n64), .S(OP2[24]), .Z(n410) );
  INV_X1 U639 ( .A(OP1[24]), .ZN(n625) );
  AOI21_X1 U640 ( .B1(n615), .B2(n410), .A(n625), .ZN(n411) );
  AOI221_X1 U641 ( .B1(OP2[24]), .B2(n413), .C1(n412), .C2(n71), .A(n411), 
        .ZN(n418) );
  AOI22_X1 U642 ( .A1(N147), .A2(n66), .B1(N180), .B2(n70), .ZN(n417) );
  NAND2_X1 U643 ( .A1(n418), .A2(n417), .ZN(RES[24]) );
  OAI21_X1 U644 ( .B1(OP1[25]), .B2(n101), .A(n98), .ZN(n422) );
  OAI211_X1 U645 ( .C1(n157), .C2(n331), .A(n356), .B(n357), .ZN(n421) );
  MUX2_X1 U646 ( .A(n101), .B(n64), .S(OP2[25]), .Z(n419) );
  INV_X1 U647 ( .A(OP1[25]), .ZN(n624) );
  AOI21_X1 U648 ( .B1(n615), .B2(n419), .A(n624), .ZN(n420) );
  AOI221_X1 U649 ( .B1(OP2[25]), .B2(n422), .C1(n421), .C2(n71), .A(n420), 
        .ZN(n428) );
  AOI22_X1 U650 ( .A1(N148), .A2(n66), .B1(N181), .B2(n70), .ZN(n427) );
  NAND2_X1 U651 ( .A1(n428), .A2(n427), .ZN(RES[25]) );
  OAI21_X1 U652 ( .B1(OP1[26]), .B2(n101), .A(n98), .ZN(n441) );
  OAI211_X1 U653 ( .C1(n344), .C2(n331), .A(n345), .B(n346), .ZN(n431) );
  MUX2_X1 U654 ( .A(n101), .B(n64), .S(n15), .Z(n429) );
  INV_X1 U655 ( .A(OP1[26]), .ZN(n623) );
  AOI21_X1 U656 ( .B1(n615), .B2(n429), .A(n623), .ZN(n430) );
  AOI221_X1 U657 ( .B1(n15), .B2(n441), .C1(n431), .C2(n71), .A(n430), .ZN(
        n443) );
  AOI22_X1 U658 ( .A1(N149), .A2(n66), .B1(N182), .B2(n70), .ZN(n442) );
  NAND2_X1 U659 ( .A1(n443), .A2(n442), .ZN(RES[26]) );
  OAI21_X1 U660 ( .B1(OP1[27]), .B2(n101), .A(n98), .ZN(n451) );
  OAI211_X1 U661 ( .C1(n261), .C2(n236), .A(n325), .B(n326), .ZN(n450) );
  MUX2_X1 U662 ( .A(n101), .B(n64), .S(OP2[27]), .Z(n444) );
  INV_X1 U663 ( .A(OP1[27]), .ZN(n622) );
  AOI21_X1 U664 ( .B1(n615), .B2(n444), .A(n622), .ZN(n445) );
  AOI221_X1 U665 ( .B1(OP2[27]), .B2(n451), .C1(n450), .C2(n71), .A(n445), 
        .ZN(n453) );
  AOI22_X1 U666 ( .A1(N150), .A2(n66), .B1(N183), .B2(n70), .ZN(n452) );
  NAND2_X1 U667 ( .A1(n452), .A2(n453), .ZN(RES[27]) );
  NAND2_X1 U668 ( .A1(n73), .A2(n6), .ZN(n495) );
  INV_X1 U669 ( .A(OP1[28]), .ZN(n621) );
  AOI21_X1 U670 ( .B1(n56), .B2(n621), .A(n99), .ZN(n455) );
  INV_X1 U671 ( .A(OP2[28]), .ZN(n454) );
  OAI22_X1 U672 ( .A1(n312), .A2(n495), .B1(n455), .B2(n454), .ZN(n461) );
  AOI21_X1 U673 ( .B1(n55), .B2(n378), .A(n461), .ZN(n465) );
  MUX2_X1 U674 ( .A(n101), .B(n64), .S(OP2[28]), .Z(n462) );
  AOI21_X1 U675 ( .B1(n615), .B2(n462), .A(n621), .ZN(n463) );
  AOI221_X1 U676 ( .B1(N184), .B2(n68), .C1(N151), .C2(n66), .A(n463), .ZN(
        n464) );
  NAND2_X1 U677 ( .A1(n465), .A2(n464), .ZN(RES[28]) );
  INV_X1 U678 ( .A(OP1[29]), .ZN(n620) );
  AOI21_X1 U679 ( .B1(n56), .B2(n620), .A(n99), .ZN(n471) );
  INV_X1 U680 ( .A(OP2[29]), .ZN(n466) );
  OAI22_X1 U681 ( .A1(n298), .A2(n495), .B1(n471), .B2(n466), .ZN(n472) );
  AOI21_X1 U682 ( .B1(n55), .B2(n363), .A(n472), .ZN(n476) );
  MUX2_X1 U683 ( .A(n101), .B(n64), .S(OP2[29]), .Z(n473) );
  AOI21_X1 U684 ( .B1(n615), .B2(n473), .A(n620), .ZN(n474) );
  AOI221_X1 U685 ( .B1(N185), .B2(n68), .C1(N152), .C2(n66), .A(n474), .ZN(
        n475) );
  NAND2_X1 U686 ( .A1(n476), .A2(n475), .ZN(RES[29]) );
  INV_X1 U687 ( .A(OP1[30]), .ZN(n619) );
  AOI21_X1 U688 ( .B1(n56), .B2(n619), .A(n99), .ZN(n482) );
  INV_X1 U689 ( .A(OP2[30]), .ZN(n481) );
  OAI22_X1 U690 ( .A1(n271), .A2(n495), .B1(n482), .B2(n481), .ZN(n483) );
  MUX2_X1 U691 ( .A(n101), .B(n64), .S(OP2[30]), .Z(n484) );
  AOI21_X1 U692 ( .B1(n615), .B2(n484), .A(n619), .ZN(n485) );
  AOI221_X1 U693 ( .B1(N186), .B2(n68), .C1(N153), .C2(n66), .A(n485), .ZN(
        n486) );
  NAND2_X1 U694 ( .A1(n486), .A2(n492), .ZN(RES[30]) );
  INV_X1 U695 ( .A(OP1[31]), .ZN(n618) );
  AOI21_X1 U696 ( .B1(n56), .B2(n618), .A(n99), .ZN(n494) );
  INV_X1 U697 ( .A(OP2[31]), .ZN(n493) );
  OAI22_X1 U698 ( .A1(n252), .A2(n495), .B1(n494), .B2(n493), .ZN(n496) );
  AOI21_X1 U699 ( .B1(n55), .B2(n5), .A(n496), .ZN(n504) );
  MUX2_X1 U700 ( .A(n101), .B(n64), .S(OP2[31]), .Z(n497) );
  AOI21_X1 U701 ( .B1(n615), .B2(n497), .A(n618), .ZN(n502) );
  NAND2_X1 U702 ( .A1(n503), .A2(n504), .ZN(RES[31]) );
  INV_X1 U703 ( .A(n378), .ZN(n649) );
  INV_X1 U704 ( .A(n235), .ZN(n710) );
  INV_X1 U705 ( .A(n363), .ZN(n641) );
  INV_X1 U706 ( .A(n405), .ZN(n645) );
  INV_X1 U707 ( .A(RES[10]), .ZN(n507) );
  INV_X1 U708 ( .A(RES[11]), .ZN(n506) );
  INV_X1 U709 ( .A(RES[1]), .ZN(n505) );
  NAND4_X1 U710 ( .A1(n507), .A2(n506), .A3(n49), .A4(n505), .ZN(n566) );
  INV_X1 U711 ( .A(RES[14]), .ZN(n521) );
  INV_X1 U712 ( .A(RES[15]), .ZN(n520) );
  INV_X1 U713 ( .A(RES[12]), .ZN(n519) );
  INV_X1 U714 ( .A(RES[13]), .ZN(n518) );
  NAND4_X1 U715 ( .A1(n521), .A2(n520), .A3(n519), .A4(n518), .ZN(n564) );
  INV_X1 U716 ( .A(RES[18]), .ZN(n531) );
  INV_X1 U717 ( .A(RES[19]), .ZN(n530) );
  INV_X1 U718 ( .A(RES[16]), .ZN(n523) );
  INV_X1 U719 ( .A(RES[17]), .ZN(n522) );
  NAND4_X1 U720 ( .A1(n531), .A2(n530), .A3(n523), .A4(n522), .ZN(n563) );
  INV_X1 U721 ( .A(RES[22]), .ZN(n549) );
  INV_X1 U722 ( .A(RES[20]), .ZN(n533) );
  INV_X1 U723 ( .A(RES[21]), .ZN(n532) );
  NAND4_X1 U724 ( .A1(n549), .A2(n548), .A3(n533), .A4(n532), .ZN(n550) );
  NOR4_X1 U725 ( .A1(n566), .A2(n564), .A3(n563), .A4(n550), .ZN(n127) );
  INV_X1 U726 ( .A(RES[4]), .ZN(n570) );
  INV_X1 U727 ( .A(RES[5]), .ZN(n569) );
  INV_X1 U728 ( .A(RES[2]), .ZN(n568) );
  INV_X1 U729 ( .A(RES[3]), .ZN(n567) );
  NAND4_X1 U730 ( .A1(n570), .A2(n569), .A3(n568), .A4(n567), .ZN(n614) );
  INV_X1 U731 ( .A(RES[8]), .ZN(n602) );
  INV_X1 U732 ( .A(RES[9]), .ZN(n575) );
  INV_X1 U733 ( .A(RES[6]), .ZN(n572) );
  INV_X1 U734 ( .A(RES[7]), .ZN(n571) );
  NAND4_X1 U735 ( .A1(n602), .A2(n575), .A3(n572), .A4(n571), .ZN(n613) );
  INV_X1 U736 ( .A(RES[26]), .ZN(n606) );
  INV_X1 U737 ( .A(RES[27]), .ZN(n605) );
  INV_X1 U738 ( .A(RES[24]), .ZN(n604) );
  INV_X1 U739 ( .A(RES[25]), .ZN(n603) );
  NAND4_X1 U740 ( .A1(n606), .A2(n605), .A3(n604), .A4(n603), .ZN(n612) );
  INV_X1 U741 ( .A(n34), .ZN(n610) );
  INV_X1 U742 ( .A(n37), .ZN(n609) );
  INV_X1 U743 ( .A(RES[28]), .ZN(n608) );
  INV_X1 U744 ( .A(RES[29]), .ZN(n607) );
  NAND4_X1 U745 ( .A1(n610), .A2(n609), .A3(n608), .A4(n607), .ZN(n611) );
  NOR4_X1 U746 ( .A1(n614), .A2(n613), .A3(n612), .A4(n611), .ZN(n128) );
endmodule


module MUX21_NBIT32_4 ( IN0, IN1, S, O );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66;

  INV_X1 U1 ( .A(n9), .ZN(n3) );
  INV_X1 U2 ( .A(n9), .ZN(n4) );
  INV_X1 U3 ( .A(n64), .ZN(O[29]) );
  AOI22_X1 U4 ( .A1(IN0[29]), .A2(n8), .B1(IN1[29]), .B2(n3), .ZN(n64) );
  INV_X1 U5 ( .A(n63), .ZN(O[28]) );
  AOI22_X1 U6 ( .A1(IN0[28]), .A2(n7), .B1(IN1[28]), .B2(n3), .ZN(n63) );
  INV_X1 U7 ( .A(n57), .ZN(O[22]) );
  AOI22_X1 U8 ( .A1(IN0[22]), .A2(n6), .B1(IN1[22]), .B2(n3), .ZN(n57) );
  INV_X1 U9 ( .A(n55), .ZN(O[20]) );
  AOI22_X1 U10 ( .A1(IN0[20]), .A2(n5), .B1(IN1[20]), .B2(n3), .ZN(n55) );
  INV_X1 U11 ( .A(n58), .ZN(O[23]) );
  AOI22_X1 U12 ( .A1(IN0[23]), .A2(n6), .B1(IN1[23]), .B2(n3), .ZN(n58) );
  INV_X1 U13 ( .A(n56), .ZN(O[21]) );
  AOI22_X1 U14 ( .A1(IN0[21]), .A2(n6), .B1(IN1[21]), .B2(n3), .ZN(n56) );
  INV_X1 U15 ( .A(n54), .ZN(O[19]) );
  AOI22_X1 U16 ( .A1(IN0[19]), .A2(n5), .B1(IN1[19]), .B2(n4), .ZN(n54) );
  INV_X1 U17 ( .A(n62), .ZN(O[27]) );
  AOI22_X1 U18 ( .A1(IN0[27]), .A2(n7), .B1(IN1[27]), .B2(n3), .ZN(n62) );
  INV_X1 U19 ( .A(n59), .ZN(O[24]) );
  AOI22_X1 U20 ( .A1(IN0[24]), .A2(n5), .B1(IN1[24]), .B2(n3), .ZN(n59) );
  INV_X1 U21 ( .A(n60), .ZN(O[25]) );
  AOI22_X1 U22 ( .A1(IN0[25]), .A2(n7), .B1(IN1[25]), .B2(n3), .ZN(n60) );
  INV_X1 U23 ( .A(n65), .ZN(O[30]) );
  AOI22_X1 U24 ( .A1(IN0[30]), .A2(n8), .B1(IN1[30]), .B2(n3), .ZN(n65) );
  INV_X1 U25 ( .A(n61), .ZN(O[26]) );
  AOI22_X1 U26 ( .A1(IN0[26]), .A2(n8), .B1(IN1[26]), .B2(n3), .ZN(n61) );
  INV_X1 U27 ( .A(n66), .ZN(O[31]) );
  AOI22_X1 U28 ( .A1(IN0[31]), .A2(n8), .B1(IN1[31]), .B2(n3), .ZN(n66) );
  CLKBUF_X1 U29 ( .A(S), .Z(n1) );
  CLKBUF_X1 U30 ( .A(S), .Z(n2) );
  INV_X1 U31 ( .A(n1), .ZN(n5) );
  INV_X1 U32 ( .A(n1), .ZN(n6) );
  INV_X1 U33 ( .A(n2), .ZN(n7) );
  INV_X1 U34 ( .A(n2), .ZN(n8) );
  INV_X1 U35 ( .A(S), .ZN(n9) );
  MUX2_X1 U36 ( .A(IN0[0]), .B(IN1[0]), .S(S), .Z(O[0]) );
  MUX2_X1 U37 ( .A(IN0[1]), .B(IN1[1]), .S(S), .Z(O[1]) );
  MUX2_X1 U38 ( .A(IN0[2]), .B(IN1[2]), .S(n4), .Z(O[2]) );
  MUX2_X1 U39 ( .A(IN0[3]), .B(IN1[3]), .S(n4), .Z(O[3]) );
  MUX2_X1 U40 ( .A(IN0[4]), .B(IN1[4]), .S(n4), .Z(O[4]) );
  MUX2_X1 U41 ( .A(IN0[5]), .B(IN1[5]), .S(n4), .Z(O[5]) );
  MUX2_X1 U42 ( .A(IN0[6]), .B(IN1[6]), .S(n4), .Z(O[6]) );
  MUX2_X1 U43 ( .A(IN0[7]), .B(IN1[7]), .S(n4), .Z(O[7]) );
  MUX2_X1 U44 ( .A(IN0[8]), .B(IN1[8]), .S(n4), .Z(O[8]) );
  MUX2_X1 U45 ( .A(IN0[9]), .B(IN1[9]), .S(n4), .Z(O[9]) );
  MUX2_X1 U46 ( .A(IN0[10]), .B(IN1[10]), .S(n4), .Z(O[10]) );
  MUX2_X1 U47 ( .A(IN0[11]), .B(IN1[11]), .S(n4), .Z(O[11]) );
  MUX2_X1 U48 ( .A(IN0[12]), .B(IN1[12]), .S(n4), .Z(O[12]) );
  MUX2_X1 U49 ( .A(IN0[13]), .B(IN1[13]), .S(n4), .Z(O[13]) );
  MUX2_X1 U50 ( .A(IN0[14]), .B(IN1[14]), .S(n4), .Z(O[14]) );
  MUX2_X1 U51 ( .A(IN0[15]), .B(IN1[15]), .S(n4), .Z(O[15]) );
  MUX2_X1 U52 ( .A(IN0[16]), .B(IN1[16]), .S(n4), .Z(O[16]) );
  MUX2_X1 U53 ( .A(IN0[17]), .B(IN1[17]), .S(n4), .Z(O[17]) );
  MUX2_X1 U54 ( .A(IN0[18]), .B(IN1[18]), .S(n4), .Z(O[18]) );
endmodule


module ADDER_1_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212;

  AND2_X1 U2 ( .A1(n12), .A2(n15), .ZN(n1) );
  XOR2_X1 U3 ( .A(n2), .B(n52), .Z(SUM[29]) );
  NAND2_X1 U4 ( .A1(n53), .A2(n54), .ZN(n2) );
  XNOR2_X1 U5 ( .A(n45), .B(n3), .ZN(SUM[31]) );
  XOR2_X1 U6 ( .A(B[31]), .B(A[31]), .Z(n3) );
  AND2_X1 U7 ( .A1(n133), .A2(n205), .ZN(SUM[0]) );
  OAI21_X1 U8 ( .B1(n204), .B2(n168), .A(n198), .ZN(n14) );
  OAI21_X1 U9 ( .B1(n181), .B2(n167), .A(n149), .ZN(n179) );
  INV_X1 U10 ( .A(n204), .ZN(n34) );
  NAND2_X1 U11 ( .A1(n151), .A2(n153), .ZN(n147) );
  OAI21_X1 U12 ( .B1(n175), .B2(n161), .A(n163), .ZN(n172) );
  OAI21_X1 U13 ( .B1(n26), .B2(n27), .A(n28), .ZN(n22) );
  OAI21_X1 U14 ( .B1(n195), .B2(n196), .A(n12), .ZN(n193) );
  OAI21_X1 U15 ( .B1(n116), .B2(n117), .A(n118), .ZN(n113) );
  NOR2_X1 U16 ( .A1(n119), .A2(n120), .ZN(n118) );
  OAI21_X1 U17 ( .B1(n91), .B2(n92), .A(n93), .ZN(n88) );
  NOR2_X1 U18 ( .A1(n7), .A2(n94), .ZN(n93) );
  AOI21_X1 U19 ( .B1(n95), .B2(n96), .A(n97), .ZN(n94) );
  OAI21_X1 U20 ( .B1(n66), .B2(n67), .A(n68), .ZN(n63) );
  NOR2_X1 U21 ( .A1(n8), .A2(n69), .ZN(n68) );
  AOI21_X1 U22 ( .B1(n70), .B2(n71), .A(n72), .ZN(n69) );
  AOI21_X1 U23 ( .B1(n121), .B2(n122), .A(n123), .ZN(n120) );
  NAND2_X1 U24 ( .A1(n125), .A2(n126), .ZN(n121) );
  OAI21_X1 U25 ( .B1(n127), .B2(n128), .A(n129), .ZN(n126) );
  NAND4_X1 U26 ( .A1(n35), .A2(n29), .A3(n21), .A4(n23), .ZN(n168) );
  NAND4_X1 U27 ( .A1(n182), .A2(n188), .A3(n11), .A4(n16), .ZN(n167) );
  OAI21_X1 U28 ( .B1(n51), .B2(n52), .A(n53), .ZN(n46) );
  AOI21_X1 U29 ( .B1(n158), .B2(n159), .A(n160), .ZN(n155) );
  OAI21_X1 U30 ( .B1(n161), .B2(n162), .A(n163), .ZN(n159) );
  AOI21_X1 U31 ( .B1(n182), .B2(n183), .A(n184), .ZN(n149) );
  INV_X1 U32 ( .A(n185), .ZN(n184) );
  OAI21_X1 U33 ( .B1(n1), .B2(n186), .A(n187), .ZN(n183) );
  NAND2_X1 U34 ( .A1(n101), .A2(n114), .ZN(n115) );
  NAND2_X1 U35 ( .A1(n185), .A2(n182), .ZN(n189) );
  NAND2_X1 U36 ( .A1(n131), .A2(n124), .ZN(n134) );
  NAND2_X1 U37 ( .A1(n43), .A2(n44), .ZN(n37) );
  NAND2_X1 U38 ( .A1(n206), .A2(n207), .ZN(n152) );
  AOI21_X1 U39 ( .B1(n209), .B2(n43), .A(n210), .ZN(n206) );
  NAND4_X1 U40 ( .A1(n208), .A2(n58), .A3(n60), .A4(n43), .ZN(n207) );
  NAND2_X1 U41 ( .A1(n116), .A2(n128), .ZN(n141) );
  NAND2_X1 U42 ( .A1(n66), .A2(n76), .ZN(n86) );
  NAND2_X1 U43 ( .A1(n91), .A2(n101), .ZN(n111) );
  NAND2_X1 U44 ( .A1(n110), .A2(n102), .ZN(n107) );
  NAND2_X1 U45 ( .A1(n103), .A2(n111), .ZN(n110) );
  NAND2_X1 U46 ( .A1(n85), .A2(n77), .ZN(n82) );
  NAND2_X1 U47 ( .A1(n78), .A2(n86), .ZN(n85) );
  OR2_X1 U48 ( .A1(n154), .A2(n5), .ZN(n143) );
  AND2_X1 U49 ( .A1(n6), .A2(n146), .ZN(n5) );
  OAI21_X1 U50 ( .B1(n155), .B2(n156), .A(n157), .ZN(n154) );
  XNOR2_X1 U51 ( .A(n107), .B(n109), .ZN(SUM[22]) );
  NAND2_X1 U52 ( .A1(n96), .A2(n98), .ZN(n109) );
  XNOR2_X1 U53 ( .A(n82), .B(n84), .ZN(SUM[26]) );
  NAND2_X1 U54 ( .A1(n71), .A2(n73), .ZN(n84) );
  XNOR2_X1 U55 ( .A(n169), .B(n170), .ZN(SUM[15]) );
  NOR2_X1 U56 ( .A1(n156), .A2(n171), .ZN(n170) );
  AOI21_X1 U57 ( .B1(n158), .B2(n172), .A(n160), .ZN(n169) );
  XNOR2_X1 U58 ( .A(n143), .B(n145), .ZN(SUM[16]) );
  NAND2_X1 U59 ( .A1(n128), .A2(n144), .ZN(n145) );
  XNOR2_X1 U60 ( .A(n17), .B(n18), .ZN(SUM[7]) );
  NAND2_X1 U61 ( .A1(n23), .A2(n24), .ZN(n17) );
  NAND2_X1 U62 ( .A1(n19), .A2(n20), .ZN(n18) );
  NAND2_X1 U63 ( .A1(n21), .A2(n22), .ZN(n19) );
  XNOR2_X1 U64 ( .A(n25), .B(n22), .ZN(SUM[6]) );
  NAND2_X1 U65 ( .A1(n21), .A2(n20), .ZN(n25) );
  XNOR2_X1 U66 ( .A(n105), .B(n106), .ZN(SUM[23]) );
  NOR2_X1 U67 ( .A1(n97), .A2(n7), .ZN(n106) );
  AOI21_X1 U68 ( .B1(n98), .B2(n107), .A(n108), .ZN(n105) );
  XNOR2_X1 U69 ( .A(n80), .B(n81), .ZN(SUM[27]) );
  NOR2_X1 U70 ( .A1(n72), .A2(n8), .ZN(n81) );
  AOI21_X1 U71 ( .B1(n73), .B2(n82), .A(n83), .ZN(n80) );
  XNOR2_X1 U72 ( .A(n9), .B(n10), .ZN(SUM[9]) );
  NAND2_X1 U73 ( .A1(n11), .A2(n12), .ZN(n9) );
  XNOR2_X1 U74 ( .A(n31), .B(n30), .ZN(SUM[5]) );
  NAND2_X1 U75 ( .A1(n29), .A2(n28), .ZN(n31) );
  XNOR2_X1 U76 ( .A(n88), .B(n90), .ZN(SUM[24]) );
  NAND2_X1 U77 ( .A1(n76), .A2(n89), .ZN(n90) );
  XNOR2_X1 U78 ( .A(n63), .B(n65), .ZN(SUM[28]) );
  NAND2_X1 U79 ( .A1(n62), .A2(n64), .ZN(n65) );
  XNOR2_X1 U80 ( .A(n36), .B(n34), .ZN(SUM[4]) );
  NAND2_X1 U81 ( .A1(n33), .A2(n35), .ZN(n36) );
  XNOR2_X1 U82 ( .A(n13), .B(n14), .ZN(SUM[8]) );
  NAND2_X1 U83 ( .A1(n15), .A2(n16), .ZN(n13) );
  XNOR2_X1 U84 ( .A(n180), .B(n179), .ZN(SUM[12]) );
  NAND2_X1 U85 ( .A1(n162), .A2(n164), .ZN(n180) );
  XNOR2_X1 U86 ( .A(n112), .B(n111), .ZN(SUM[21]) );
  NAND2_X1 U87 ( .A1(n102), .A2(n103), .ZN(n112) );
  XNOR2_X1 U88 ( .A(n87), .B(n86), .ZN(SUM[25]) );
  NAND2_X1 U89 ( .A1(n77), .A2(n78), .ZN(n87) );
  XNOR2_X1 U90 ( .A(n142), .B(n141), .ZN(SUM[17]) );
  NAND2_X1 U91 ( .A1(n129), .A2(n130), .ZN(n142) );
  XNOR2_X1 U92 ( .A(n177), .B(n176), .ZN(SUM[13]) );
  NAND2_X1 U93 ( .A1(n163), .A2(n165), .ZN(n177) );
  XNOR2_X1 U94 ( .A(n132), .B(n59), .ZN(SUM[1]) );
  NAND2_X1 U95 ( .A1(n58), .A2(n57), .ZN(n132) );
  XNOR2_X1 U96 ( .A(n139), .B(n138), .ZN(SUM[18]) );
  NAND2_X1 U97 ( .A1(n122), .A2(n125), .ZN(n139) );
  XNOR2_X1 U98 ( .A(n55), .B(n42), .ZN(SUM[2]) );
  NAND2_X1 U99 ( .A1(n60), .A2(n41), .ZN(n55) );
  XNOR2_X1 U100 ( .A(n194), .B(n193), .ZN(SUM[10]) );
  NAND2_X1 U101 ( .A1(n187), .A2(n188), .ZN(n194) );
  XNOR2_X1 U102 ( .A(n46), .B(n50), .ZN(SUM[30]) );
  NAND2_X1 U103 ( .A1(n49), .A2(n47), .ZN(n50) );
  XNOR2_X1 U104 ( .A(n174), .B(n172), .ZN(SUM[14]) );
  NAND2_X1 U105 ( .A1(n173), .A2(n158), .ZN(n174) );
  NAND2_X1 U106 ( .A1(n197), .A2(n15), .ZN(n10) );
  NAND2_X1 U107 ( .A1(n14), .A2(n16), .ZN(n197) );
  NAND2_X1 U108 ( .A1(n32), .A2(n33), .ZN(n30) );
  NAND2_X1 U109 ( .A1(n34), .A2(n35), .ZN(n32) );
  NAND2_X1 U110 ( .A1(n178), .A2(n162), .ZN(n176) );
  NAND2_X1 U111 ( .A1(n179), .A2(n164), .ZN(n178) );
  NAND2_X1 U112 ( .A1(n140), .A2(n129), .ZN(n138) );
  NAND2_X1 U113 ( .A1(n130), .A2(n141), .ZN(n140) );
  INV_X1 U114 ( .A(n133), .ZN(n59) );
  NAND2_X1 U115 ( .A1(n143), .A2(n144), .ZN(n116) );
  NAND2_X1 U116 ( .A1(n88), .A2(n89), .ZN(n66) );
  NAND2_X1 U117 ( .A1(n113), .A2(n114), .ZN(n91) );
  NAND2_X1 U118 ( .A1(n199), .A2(n200), .ZN(n153) );
  AOI21_X1 U119 ( .B1(n202), .B2(n23), .A(n203), .ZN(n199) );
  NAND4_X1 U120 ( .A1(n201), .A2(n29), .A3(n21), .A4(n23), .ZN(n200) );
  AND2_X1 U121 ( .A1(n61), .A2(n62), .ZN(n52) );
  NAND2_X1 U122 ( .A1(n63), .A2(n64), .ZN(n61) );
  NAND2_X1 U123 ( .A1(n188), .A2(n11), .ZN(n186) );
  NAND2_X1 U124 ( .A1(n28), .A2(n33), .ZN(n201) );
  NAND2_X1 U125 ( .A1(n57), .A2(n133), .ZN(n208) );
  NAND2_X1 U126 ( .A1(n98), .A2(n99), .ZN(n95) );
  OAI21_X1 U127 ( .B1(n100), .B2(n101), .A(n102), .ZN(n99) );
  NAND2_X1 U128 ( .A1(n73), .A2(n74), .ZN(n70) );
  OAI21_X1 U129 ( .B1(n75), .B2(n76), .A(n77), .ZN(n74) );
  NAND2_X1 U130 ( .A1(n56), .A2(n57), .ZN(n42) );
  NAND2_X1 U131 ( .A1(n58), .A2(n59), .ZN(n56) );
  AND4_X1 U132 ( .A1(n164), .A2(n165), .A3(n158), .A4(n166), .ZN(n6) );
  INV_X1 U133 ( .A(B[0]), .ZN(n211) );
  OR2_X1 U134 ( .A1(B[7]), .A2(A[7]), .ZN(n23) );
  OR2_X1 U135 ( .A1(B[14]), .A2(A[14]), .ZN(n158) );
  OR2_X1 U136 ( .A1(B[6]), .A2(A[6]), .ZN(n21) );
  OR2_X1 U137 ( .A1(B[9]), .A2(A[9]), .ZN(n11) );
  OR2_X1 U138 ( .A1(B[10]), .A2(A[10]), .ZN(n188) );
  OR2_X1 U139 ( .A1(B[22]), .A2(A[22]), .ZN(n98) );
  AND2_X1 U140 ( .A1(B[23]), .A2(A[23]), .ZN(n7) );
  AND2_X1 U141 ( .A1(B[27]), .A2(A[27]), .ZN(n8) );
  OR2_X1 U142 ( .A1(B[8]), .A2(A[8]), .ZN(n16) );
  OR2_X1 U143 ( .A1(B[3]), .A2(A[3]), .ZN(n43) );
  OR2_X1 U144 ( .A1(B[17]), .A2(A[17]), .ZN(n130) );
  OR2_X1 U145 ( .A1(B[21]), .A2(A[21]), .ZN(n103) );
  NAND2_X1 U146 ( .A1(B[1]), .A2(A[1]), .ZN(n57) );
  NAND2_X1 U147 ( .A1(B[8]), .A2(A[8]), .ZN(n15) );
  NAND2_X1 U148 ( .A1(B[4]), .A2(A[4]), .ZN(n33) );
  NAND2_X1 U149 ( .A1(B[16]), .A2(A[16]), .ZN(n128) );
  NAND2_X1 U150 ( .A1(B[20]), .A2(A[20]), .ZN(n101) );
  NAND2_X1 U151 ( .A1(B[12]), .A2(A[12]), .ZN(n162) );
  NAND2_X1 U152 ( .A1(B[24]), .A2(A[24]), .ZN(n76) );
  OR2_X1 U153 ( .A1(B[12]), .A2(A[12]), .ZN(n164) );
  OR2_X1 U154 ( .A1(B[4]), .A2(A[4]), .ZN(n35) );
  NAND2_X1 U155 ( .A1(B[0]), .A2(A[0]), .ZN(n133) );
  NAND2_X1 U156 ( .A1(B[17]), .A2(A[17]), .ZN(n129) );
  NAND2_X1 U157 ( .A1(B[21]), .A2(A[21]), .ZN(n102) );
  NAND2_X1 U158 ( .A1(B[9]), .A2(A[9]), .ZN(n12) );
  NAND2_X1 U159 ( .A1(B[5]), .A2(A[5]), .ZN(n28) );
  NAND2_X1 U160 ( .A1(B[25]), .A2(A[25]), .ZN(n77) );
  OR2_X1 U161 ( .A1(B[11]), .A2(A[11]), .ZN(n182) );
  NAND2_X1 U162 ( .A1(B[13]), .A2(A[13]), .ZN(n163) );
  OR2_X1 U163 ( .A1(B[1]), .A2(A[1]), .ZN(n58) );
  NAND2_X1 U164 ( .A1(B[6]), .A2(A[6]), .ZN(n20) );
  OR2_X1 U165 ( .A1(B[13]), .A2(A[13]), .ZN(n165) );
  NAND2_X1 U166 ( .A1(B[22]), .A2(A[22]), .ZN(n96) );
  NAND2_X1 U167 ( .A1(B[26]), .A2(A[26]), .ZN(n71) );
  NAND2_X1 U168 ( .A1(B[18]), .A2(A[18]), .ZN(n122) );
  OR2_X1 U169 ( .A1(B[2]), .A2(A[2]), .ZN(n60) );
  NAND2_X1 U170 ( .A1(B[10]), .A2(A[10]), .ZN(n187) );
  NAND2_X1 U171 ( .A1(B[2]), .A2(A[2]), .ZN(n41) );
  OR2_X1 U172 ( .A1(B[19]), .A2(A[19]), .ZN(n124) );
  OR2_X1 U173 ( .A1(B[16]), .A2(A[16]), .ZN(n144) );
  OR2_X1 U174 ( .A1(B[20]), .A2(A[20]), .ZN(n114) );
  OR2_X1 U175 ( .A1(B[24]), .A2(A[24]), .ZN(n89) );
  NAND2_X1 U176 ( .A1(B[11]), .A2(A[11]), .ZN(n185) );
  NAND2_X1 U177 ( .A1(B[29]), .A2(A[29]), .ZN(n53) );
  OR2_X1 U178 ( .A1(B[15]), .A2(A[15]), .ZN(n166) );
  NAND2_X1 U179 ( .A1(B[3]), .A2(A[3]), .ZN(n44) );
  NAND2_X1 U180 ( .A1(B[7]), .A2(A[7]), .ZN(n24) );
  NAND2_X1 U181 ( .A1(B[15]), .A2(A[15]), .ZN(n157) );
  OR2_X1 U182 ( .A1(B[29]), .A2(A[29]), .ZN(n54) );
  OR2_X1 U183 ( .A1(B[30]), .A2(A[30]), .ZN(n47) );
  NAND2_X1 U184 ( .A1(B[28]), .A2(A[28]), .ZN(n62) );
  NAND2_X1 U185 ( .A1(B[14]), .A2(A[14]), .ZN(n173) );
  NAND2_X1 U186 ( .A1(B[19]), .A2(A[19]), .ZN(n131) );
  NAND2_X1 U187 ( .A1(B[30]), .A2(A[30]), .ZN(n49) );
  OR2_X1 U188 ( .A1(B[27]), .A2(A[27]), .ZN(n79) );
  OR2_X1 U189 ( .A1(B[18]), .A2(A[18]), .ZN(n125) );
  OR2_X1 U190 ( .A1(B[5]), .A2(A[5]), .ZN(n29) );
  OR2_X1 U191 ( .A1(B[23]), .A2(A[23]), .ZN(n104) );
  OR2_X1 U192 ( .A1(B[28]), .A2(A[28]), .ZN(n64) );
  OR2_X1 U193 ( .A1(B[25]), .A2(A[25]), .ZN(n78) );
  OR2_X1 U194 ( .A1(B[26]), .A2(A[26]), .ZN(n73) );
  NAND2_X1 U195 ( .A1(n211), .A2(n212), .ZN(n205) );
  INV_X1 U196 ( .A(A[0]), .ZN(n212) );
  INV_X1 U197 ( .A(n29), .ZN(n27) );
  INV_X1 U198 ( .A(n30), .ZN(n26) );
  XNOR2_X1 U199 ( .A(n37), .B(n38), .ZN(SUM[3]) );
  OAI21_X1 U200 ( .B1(n39), .B2(n40), .A(n41), .ZN(n38) );
  INV_X1 U201 ( .A(n42), .ZN(n39) );
  AOI21_X1 U202 ( .B1(n46), .B2(n47), .A(n48), .ZN(n45) );
  INV_X1 U203 ( .A(n49), .ZN(n48) );
  INV_X1 U204 ( .A(n54), .ZN(n51) );
  INV_X1 U205 ( .A(n78), .ZN(n75) );
  NAND3_X1 U206 ( .A1(n73), .A2(n79), .A3(n78), .ZN(n67) );
  INV_X1 U207 ( .A(n79), .ZN(n72) );
  INV_X1 U208 ( .A(n71), .ZN(n83) );
  INV_X1 U209 ( .A(n103), .ZN(n100) );
  NAND3_X1 U210 ( .A1(n98), .A2(n104), .A3(n103), .ZN(n92) );
  INV_X1 U211 ( .A(n104), .ZN(n97) );
  INV_X1 U212 ( .A(n96), .ZN(n108) );
  XNOR2_X1 U213 ( .A(n115), .B(n113), .ZN(SUM[20]) );
  INV_X1 U214 ( .A(n124), .ZN(n123) );
  INV_X1 U215 ( .A(n130), .ZN(n127) );
  INV_X1 U216 ( .A(n131), .ZN(n119) );
  NAND3_X1 U217 ( .A1(n125), .A2(n124), .A3(n130), .ZN(n117) );
  XNOR2_X1 U218 ( .A(n134), .B(n135), .ZN(SUM[19]) );
  OAI21_X1 U219 ( .B1(n136), .B2(n137), .A(n122), .ZN(n135) );
  INV_X1 U220 ( .A(n125), .ZN(n137) );
  INV_X1 U221 ( .A(n138), .ZN(n136) );
  NAND3_X1 U222 ( .A1(n147), .A2(n148), .A3(n149), .ZN(n146) );
  NAND3_X1 U223 ( .A1(n150), .A2(n151), .A3(n152), .ZN(n148) );
  INV_X1 U224 ( .A(n167), .ZN(n151) );
  INV_X1 U225 ( .A(n168), .ZN(n150) );
  INV_X1 U226 ( .A(n157), .ZN(n171) );
  INV_X1 U227 ( .A(n166), .ZN(n156) );
  INV_X1 U228 ( .A(n173), .ZN(n160) );
  INV_X1 U229 ( .A(n165), .ZN(n161) );
  INV_X1 U230 ( .A(n176), .ZN(n175) );
  INV_X1 U231 ( .A(n14), .ZN(n181) );
  XNOR2_X1 U232 ( .A(n189), .B(n190), .ZN(SUM[11]) );
  OAI21_X1 U233 ( .B1(n191), .B2(n192), .A(n187), .ZN(n190) );
  INV_X1 U234 ( .A(n188), .ZN(n192) );
  INV_X1 U235 ( .A(n193), .ZN(n191) );
  INV_X1 U236 ( .A(n10), .ZN(n196) );
  INV_X1 U237 ( .A(n153), .ZN(n198) );
  INV_X1 U238 ( .A(n24), .ZN(n203) );
  INV_X1 U239 ( .A(n20), .ZN(n202) );
  INV_X1 U240 ( .A(n60), .ZN(n40) );
  INV_X1 U241 ( .A(n152), .ZN(n204) );
  INV_X1 U242 ( .A(n44), .ZN(n210) );
  INV_X1 U243 ( .A(n41), .ZN(n209) );
  INV_X1 U244 ( .A(n11), .ZN(n195) );
endmodule


module ADDER_1 ( A, B, S );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;


  ADDER_1_DW01_add_2 add_16 ( .A(A), .B(B), .CI(1'b0), .SUM(S) );
endmodule


module MUX21_NBIT32_3 ( IN0, IN1, S, O );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  INV_X1 U3 ( .A(n94), .ZN(O[23]) );
  INV_X1 U4 ( .A(n85), .ZN(O[15]) );
  INV_X1 U5 ( .A(n103), .ZN(O[31]) );
  INV_X1 U6 ( .A(n110), .ZN(O[9]) );
  INV_X1 U7 ( .A(n109), .ZN(O[8]) );
  INV_X1 U8 ( .A(n108), .ZN(O[7]) );
  INV_X1 U9 ( .A(n107), .ZN(O[6]) );
  INV_X1 U10 ( .A(n106), .ZN(O[5]) );
  INV_X1 U11 ( .A(n105), .ZN(O[4]) );
  INV_X1 U12 ( .A(n104), .ZN(O[3]) );
  INV_X1 U13 ( .A(n86), .ZN(O[16]) );
  INV_X1 U14 ( .A(n93), .ZN(O[22]) );
  INV_X1 U15 ( .A(n100), .ZN(O[29]) );
  INV_X1 U16 ( .A(n97), .ZN(O[26]) );
  INV_X1 U17 ( .A(n96), .ZN(O[25]) );
  INV_X1 U18 ( .A(n95), .ZN(O[24]) );
  INV_X1 U19 ( .A(n92), .ZN(O[21]) );
  INV_X1 U20 ( .A(n91), .ZN(O[20]) );
  INV_X1 U21 ( .A(n84), .ZN(O[14]) );
  INV_X1 U22 ( .A(n83), .ZN(O[13]) );
  INV_X1 U23 ( .A(n82), .ZN(O[12]) );
  INV_X1 U24 ( .A(n102), .ZN(O[30]) );
  INV_X1 U25 ( .A(n99), .ZN(O[28]) );
  INV_X1 U26 ( .A(n89), .ZN(O[19]) );
  INV_X1 U27 ( .A(n88), .ZN(O[18]) );
  INV_X1 U28 ( .A(n87), .ZN(O[17]) );
  INV_X1 U29 ( .A(n81), .ZN(O[11]) );
  INV_X1 U30 ( .A(n80), .ZN(O[10]) );
  INV_X1 U31 ( .A(n101), .ZN(O[2]) );
  INV_X1 U32 ( .A(n90), .ZN(O[1]) );
  INV_X1 U33 ( .A(n79), .ZN(O[0]) );
  BUF_X1 U34 ( .A(n2), .Z(n11) );
  BUF_X1 U35 ( .A(n1), .Z(n6) );
  BUF_X1 U36 ( .A(n1), .Z(n7) );
  BUF_X1 U37 ( .A(n2), .Z(n10) );
  BUF_X1 U38 ( .A(n3), .Z(n14) );
  BUF_X1 U39 ( .A(n3), .Z(n13) );
  BUF_X1 U40 ( .A(n1), .Z(n8) );
  BUF_X1 U41 ( .A(n2), .Z(n9) );
  BUF_X1 U42 ( .A(n3), .Z(n12) );
  AOI22_X1 U43 ( .A1(IN0[31]), .A2(n4), .B1(IN1[31]), .B2(n7), .ZN(n103) );
  AOI22_X1 U44 ( .A1(IN0[9]), .A2(n5), .B1(n13), .B2(IN1[9]), .ZN(n110) );
  AOI22_X1 U45 ( .A1(IN0[8]), .A2(n4), .B1(IN1[8]), .B2(n6), .ZN(n109) );
  AOI22_X1 U46 ( .A1(IN0[7]), .A2(n5), .B1(IN1[7]), .B2(n6), .ZN(n108) );
  AOI22_X1 U47 ( .A1(IN0[6]), .A2(n4), .B1(IN1[6]), .B2(n6), .ZN(n107) );
  AOI22_X1 U48 ( .A1(IN0[5]), .A2(n5), .B1(IN1[5]), .B2(n6), .ZN(n106) );
  AOI22_X1 U49 ( .A1(IN0[4]), .A2(n4), .B1(IN1[4]), .B2(n7), .ZN(n105) );
  AOI22_X1 U50 ( .A1(IN0[3]), .A2(n5), .B1(IN1[3]), .B2(n7), .ZN(n104) );
  AOI22_X1 U51 ( .A1(IN0[30]), .A2(n5), .B1(IN1[30]), .B2(n10), .ZN(n102) );
  AOI22_X1 U52 ( .A1(IN0[29]), .A2(n5), .B1(IN1[29]), .B2(n8), .ZN(n100) );
  AOI22_X1 U53 ( .A1(IN0[28]), .A2(n5), .B1(IN1[28]), .B2(n8), .ZN(n99) );
  AOI22_X1 U54 ( .A1(IN0[26]), .A2(n5), .B1(IN1[26]), .B2(n8), .ZN(n97) );
  AOI22_X1 U55 ( .A1(IN0[25]), .A2(n5), .B1(IN1[25]), .B2(n9), .ZN(n96) );
  AOI22_X1 U56 ( .A1(IN0[24]), .A2(n5), .B1(IN1[24]), .B2(n9), .ZN(n95) );
  AOI22_X1 U57 ( .A1(IN0[22]), .A2(n5), .B1(IN1[22]), .B2(n9), .ZN(n93) );
  AOI22_X1 U58 ( .A1(IN0[21]), .A2(n5), .B1(IN1[21]), .B2(n10), .ZN(n92) );
  AOI22_X1 U59 ( .A1(IN0[20]), .A2(n5), .B1(IN1[20]), .B2(n10), .ZN(n91) );
  AOI22_X1 U60 ( .A1(IN0[19]), .A2(n4), .B1(IN1[19]), .B2(n11), .ZN(n89) );
  AOI22_X1 U61 ( .A1(IN0[18]), .A2(n4), .B1(IN1[18]), .B2(n11), .ZN(n88) );
  AOI22_X1 U62 ( .A1(IN0[17]), .A2(n4), .B1(IN1[17]), .B2(n11), .ZN(n87) );
  AOI22_X1 U63 ( .A1(IN0[16]), .A2(n4), .B1(IN1[16]), .B2(n11), .ZN(n86) );
  AOI22_X1 U64 ( .A1(IN0[14]), .A2(n4), .B1(IN1[14]), .B2(n12), .ZN(n84) );
  AOI22_X1 U65 ( .A1(IN0[13]), .A2(n4), .B1(IN1[13]), .B2(n12), .ZN(n83) );
  AOI22_X1 U66 ( .A1(IN0[12]), .A2(n4), .B1(IN1[12]), .B2(n12), .ZN(n82) );
  AOI22_X1 U67 ( .A1(IN0[11]), .A2(n4), .B1(IN1[11]), .B2(n13), .ZN(n81) );
  AOI22_X1 U68 ( .A1(IN0[10]), .A2(n4), .B1(IN1[10]), .B2(n13), .ZN(n80) );
  AOI22_X1 U69 ( .A1(IN0[2]), .A2(n5), .B1(IN1[2]), .B2(n7), .ZN(n101) );
  AOI22_X1 U70 ( .A1(IN0[1]), .A2(n4), .B1(IN1[1]), .B2(n10), .ZN(n90) );
  AOI22_X1 U71 ( .A1(IN0[0]), .A2(n4), .B1(IN1[0]), .B2(n13), .ZN(n79) );
  BUF_X1 U72 ( .A(S), .Z(n3) );
  BUF_X1 U73 ( .A(S), .Z(n1) );
  BUF_X1 U74 ( .A(S), .Z(n2) );
  INV_X1 U75 ( .A(n98), .ZN(O[27]) );
  AOI22_X1 U76 ( .A1(IN0[27]), .A2(n5), .B1(IN1[27]), .B2(n8), .ZN(n98) );
  AOI22_X1 U77 ( .A1(IN0[15]), .A2(n4), .B1(IN1[15]), .B2(n12), .ZN(n85) );
  AOI22_X1 U78 ( .A1(IN0[23]), .A2(n5), .B1(IN1[23]), .B2(n9), .ZN(n94) );
endmodule


module MUX21_NBIT32_2 ( IN0, IN1, S, O );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] O;
  input S;
  wire   n1, n2, n3, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100;

  BUF_X1 U1 ( .A(n68), .Z(n1) );
  BUF_X1 U2 ( .A(n68), .Z(n2) );
  BUF_X1 U3 ( .A(n68), .Z(n3) );
  INV_X1 U4 ( .A(n81), .ZN(O[20]) );
  INV_X1 U5 ( .A(n82), .ZN(O[21]) );
  INV_X1 U6 ( .A(n83), .ZN(O[22]) );
  INV_X1 U7 ( .A(n84), .ZN(O[23]) );
  INV_X1 U8 ( .A(n85), .ZN(O[24]) );
  INV_X1 U9 ( .A(n86), .ZN(O[25]) );
  INV_X1 U10 ( .A(n87), .ZN(O[26]) );
  INV_X1 U11 ( .A(n88), .ZN(O[27]) );
  INV_X1 U12 ( .A(n89), .ZN(O[28]) );
  INV_X1 U13 ( .A(n90), .ZN(O[29]) );
  INV_X1 U14 ( .A(n92), .ZN(O[30]) );
  INV_X1 U15 ( .A(n93), .ZN(O[31]) );
  AOI22_X1 U16 ( .A1(IN0[0]), .A2(n1), .B1(IN1[0]), .B2(S), .ZN(n69) );
  AOI22_X1 U17 ( .A1(IN0[1]), .A2(n1), .B1(IN1[1]), .B2(S), .ZN(n80) );
  AOI22_X1 U18 ( .A1(IN0[2]), .A2(n2), .B1(IN1[2]), .B2(S), .ZN(n91) );
  AOI22_X1 U19 ( .A1(IN0[3]), .A2(n3), .B1(IN1[3]), .B2(S), .ZN(n94) );
  AOI22_X1 U20 ( .A1(IN0[4]), .A2(n3), .B1(IN1[4]), .B2(S), .ZN(n95) );
  AOI22_X1 U21 ( .A1(IN0[5]), .A2(n3), .B1(IN1[5]), .B2(S), .ZN(n96) );
  AOI22_X1 U22 ( .A1(IN0[6]), .A2(n3), .B1(IN1[6]), .B2(S), .ZN(n97) );
  AOI22_X1 U23 ( .A1(IN0[7]), .A2(n3), .B1(IN1[7]), .B2(S), .ZN(n98) );
  AOI22_X1 U24 ( .A1(IN0[8]), .A2(n3), .B1(IN1[8]), .B2(S), .ZN(n99) );
  AOI22_X1 U25 ( .A1(IN0[10]), .A2(n1), .B1(IN1[10]), .B2(S), .ZN(n70) );
  AOI22_X1 U26 ( .A1(IN0[11]), .A2(n1), .B1(IN1[11]), .B2(S), .ZN(n71) );
  AOI22_X1 U27 ( .A1(IN0[12]), .A2(n1), .B1(IN1[12]), .B2(S), .ZN(n72) );
  AOI22_X1 U28 ( .A1(IN0[13]), .A2(n1), .B1(IN1[13]), .B2(S), .ZN(n73) );
  AOI22_X1 U29 ( .A1(IN0[14]), .A2(n1), .B1(IN1[14]), .B2(S), .ZN(n74) );
  AOI22_X1 U30 ( .A1(IN0[15]), .A2(n1), .B1(IN1[15]), .B2(S), .ZN(n75) );
  AOI22_X1 U31 ( .A1(IN0[16]), .A2(n1), .B1(IN1[16]), .B2(S), .ZN(n76) );
  AOI22_X1 U32 ( .A1(IN0[17]), .A2(n1), .B1(IN1[17]), .B2(S), .ZN(n77) );
  AOI22_X1 U33 ( .A1(IN0[18]), .A2(n1), .B1(IN1[18]), .B2(S), .ZN(n78) );
  AOI22_X1 U34 ( .A1(IN0[19]), .A2(n1), .B1(IN1[19]), .B2(S), .ZN(n79) );
  AOI22_X1 U35 ( .A1(IN0[20]), .A2(n2), .B1(IN1[20]), .B2(S), .ZN(n81) );
  AOI22_X1 U36 ( .A1(IN0[21]), .A2(n2), .B1(IN1[21]), .B2(S), .ZN(n82) );
  AOI22_X1 U37 ( .A1(IN0[22]), .A2(n2), .B1(IN1[22]), .B2(S), .ZN(n83) );
  AOI22_X1 U38 ( .A1(IN0[23]), .A2(n2), .B1(IN1[23]), .B2(S), .ZN(n84) );
  AOI22_X1 U39 ( .A1(IN0[24]), .A2(n2), .B1(IN1[24]), .B2(S), .ZN(n85) );
  AOI22_X1 U40 ( .A1(IN0[25]), .A2(n2), .B1(IN1[25]), .B2(S), .ZN(n86) );
  AOI22_X1 U41 ( .A1(IN0[26]), .A2(n2), .B1(IN1[26]), .B2(S), .ZN(n87) );
  AOI22_X1 U42 ( .A1(IN0[27]), .A2(n2), .B1(IN1[27]), .B2(S), .ZN(n88) );
  AOI22_X1 U43 ( .A1(IN0[28]), .A2(n2), .B1(IN1[28]), .B2(S), .ZN(n89) );
  AOI22_X1 U44 ( .A1(IN0[29]), .A2(n2), .B1(IN1[29]), .B2(S), .ZN(n90) );
  AOI22_X1 U45 ( .A1(IN0[30]), .A2(n2), .B1(IN1[30]), .B2(S), .ZN(n92) );
  AOI22_X1 U46 ( .A1(IN0[31]), .A2(n3), .B1(IN1[31]), .B2(S), .ZN(n93) );
  AOI22_X1 U47 ( .A1(IN0[9]), .A2(n3), .B1(S), .B2(IN1[9]), .ZN(n100) );
  INV_X1 U48 ( .A(n99), .ZN(O[8]) );
  INV_X1 U49 ( .A(n100), .ZN(O[9]) );
  INV_X1 U50 ( .A(n70), .ZN(O[10]) );
  INV_X1 U51 ( .A(n71), .ZN(O[11]) );
  INV_X1 U52 ( .A(n72), .ZN(O[12]) );
  INV_X1 U53 ( .A(n73), .ZN(O[13]) );
  INV_X1 U54 ( .A(n74), .ZN(O[14]) );
  INV_X1 U55 ( .A(n75), .ZN(O[15]) );
  INV_X1 U56 ( .A(n76), .ZN(O[16]) );
  INV_X1 U57 ( .A(n77), .ZN(O[17]) );
  INV_X1 U58 ( .A(n78), .ZN(O[18]) );
  INV_X1 U59 ( .A(n79), .ZN(O[19]) );
  INV_X1 U60 ( .A(n69), .ZN(O[0]) );
  INV_X1 U61 ( .A(n80), .ZN(O[1]) );
  INV_X1 U62 ( .A(n91), .ZN(O[2]) );
  INV_X1 U63 ( .A(n94), .ZN(O[3]) );
  INV_X1 U64 ( .A(n95), .ZN(O[4]) );
  INV_X1 U65 ( .A(n96), .ZN(O[5]) );
  INV_X1 U66 ( .A(n97), .ZN(O[6]) );
  INV_X1 U67 ( .A(n98), .ZN(O[7]) );
  INV_X1 U68 ( .A(S), .ZN(n68) );
endmodule


module MUX21_NBIT32_1 ( IN0, IN1, S, O );
  input [31:0] IN0;
  input [31:0] IN1;
  output [31:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n7) );
  BUF_X1 U4 ( .A(n2), .Z(n10) );
  BUF_X1 U5 ( .A(n2), .Z(n9) );
  BUF_X1 U6 ( .A(n1), .Z(n8) );
  BUF_X1 U7 ( .A(n1), .Z(n6) );
  BUF_X1 U8 ( .A(n3), .Z(n12) );
  BUF_X1 U9 ( .A(n2), .Z(n11) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(S), .Z(n3) );
  BUF_X1 U13 ( .A(S), .Z(n1) );
  BUF_X1 U14 ( .A(S), .Z(n2) );
  INV_X1 U15 ( .A(n102), .ZN(O[30]) );
  AOI22_X1 U16 ( .A1(IN0[30]), .A2(n5), .B1(IN1[30]), .B2(n10), .ZN(n102) );
  INV_X1 U17 ( .A(n81), .ZN(O[11]) );
  AOI22_X1 U18 ( .A1(IN0[11]), .A2(n4), .B1(IN1[11]), .B2(n13), .ZN(n81) );
  INV_X1 U19 ( .A(n106), .ZN(O[5]) );
  AOI22_X1 U20 ( .A1(IN0[5]), .A2(n4), .B1(IN1[5]), .B2(n6), .ZN(n106) );
  INV_X1 U21 ( .A(n80), .ZN(O[10]) );
  AOI22_X1 U22 ( .A1(IN0[10]), .A2(n4), .B1(IN1[10]), .B2(n13), .ZN(n80) );
  INV_X1 U23 ( .A(n107), .ZN(O[6]) );
  AOI22_X1 U24 ( .A1(IN0[6]), .A2(n5), .B1(IN1[6]), .B2(n6), .ZN(n107) );
  INV_X1 U25 ( .A(n108), .ZN(O[7]) );
  AOI22_X1 U26 ( .A1(IN0[7]), .A2(n4), .B1(IN1[7]), .B2(n6), .ZN(n108) );
  INV_X1 U27 ( .A(n109), .ZN(O[8]) );
  AOI22_X1 U28 ( .A1(IN0[8]), .A2(n5), .B1(IN1[8]), .B2(n6), .ZN(n109) );
  INV_X1 U29 ( .A(n110), .ZN(O[9]) );
  AOI22_X1 U30 ( .A1(IN0[9]), .A2(n4), .B1(n13), .B2(IN1[9]), .ZN(n110) );
  INV_X1 U31 ( .A(n87), .ZN(O[17]) );
  AOI22_X1 U32 ( .A1(IN0[17]), .A2(n4), .B1(IN1[17]), .B2(n11), .ZN(n87) );
  INV_X1 U33 ( .A(n82), .ZN(O[12]) );
  AOI22_X1 U34 ( .A1(IN0[12]), .A2(n4), .B1(IN1[12]), .B2(n12), .ZN(n82) );
  INV_X1 U35 ( .A(n88), .ZN(O[18]) );
  AOI22_X1 U36 ( .A1(IN0[18]), .A2(n4), .B1(IN1[18]), .B2(n11), .ZN(n88) );
  INV_X1 U37 ( .A(n86), .ZN(O[16]) );
  AOI22_X1 U38 ( .A1(IN0[16]), .A2(n4), .B1(IN1[16]), .B2(n11), .ZN(n86) );
  INV_X1 U39 ( .A(n83), .ZN(O[13]) );
  AOI22_X1 U40 ( .A1(IN0[13]), .A2(n4), .B1(IN1[13]), .B2(n12), .ZN(n83) );
  INV_X1 U41 ( .A(n85), .ZN(O[15]) );
  AOI22_X1 U42 ( .A1(IN0[15]), .A2(n4), .B1(IN1[15]), .B2(n12), .ZN(n85) );
  INV_X1 U43 ( .A(n84), .ZN(O[14]) );
  AOI22_X1 U44 ( .A1(IN0[14]), .A2(n4), .B1(IN1[14]), .B2(n12), .ZN(n84) );
  INV_X1 U45 ( .A(n104), .ZN(O[3]) );
  AOI22_X1 U46 ( .A1(IN0[3]), .A2(n5), .B1(IN1[3]), .B2(n7), .ZN(n104) );
  INV_X1 U47 ( .A(n89), .ZN(O[19]) );
  AOI22_X1 U48 ( .A1(IN0[19]), .A2(n4), .B1(IN1[19]), .B2(n11), .ZN(n89) );
  AOI22_X1 U49 ( .A1(IN0[4]), .A2(n4), .B1(IN1[4]), .B2(n7), .ZN(n105) );
  INV_X1 U50 ( .A(n90), .ZN(O[1]) );
  AOI22_X1 U51 ( .A1(IN0[1]), .A2(n4), .B1(IN1[1]), .B2(n10), .ZN(n90) );
  INV_X1 U52 ( .A(n95), .ZN(O[24]) );
  AOI22_X1 U53 ( .A1(IN0[24]), .A2(n5), .B1(IN1[24]), .B2(n9), .ZN(n95) );
  INV_X1 U54 ( .A(n94), .ZN(O[23]) );
  AOI22_X1 U55 ( .A1(IN0[23]), .A2(n5), .B1(IN1[23]), .B2(n9), .ZN(n94) );
  INV_X1 U56 ( .A(n96), .ZN(O[25]) );
  AOI22_X1 U57 ( .A1(IN0[25]), .A2(n5), .B1(IN1[25]), .B2(n9), .ZN(n96) );
  INV_X1 U58 ( .A(n97), .ZN(O[26]) );
  AOI22_X1 U59 ( .A1(IN0[26]), .A2(n5), .B1(IN1[26]), .B2(n8), .ZN(n97) );
  INV_X1 U60 ( .A(n98), .ZN(O[27]) );
  AOI22_X1 U61 ( .A1(IN0[27]), .A2(n5), .B1(IN1[27]), .B2(n8), .ZN(n98) );
  AOI22_X1 U62 ( .A1(IN0[2]), .A2(n5), .B1(IN1[2]), .B2(n7), .ZN(n101) );
  INV_X1 U63 ( .A(n91), .ZN(O[20]) );
  AOI22_X1 U64 ( .A1(IN0[20]), .A2(n5), .B1(IN1[20]), .B2(n10), .ZN(n91) );
  INV_X1 U65 ( .A(n92), .ZN(O[21]) );
  AOI22_X1 U66 ( .A1(IN0[21]), .A2(n5), .B1(IN1[21]), .B2(n10), .ZN(n92) );
  INV_X1 U67 ( .A(n93), .ZN(O[22]) );
  AOI22_X1 U68 ( .A1(IN0[22]), .A2(n5), .B1(IN1[22]), .B2(n9), .ZN(n93) );
  INV_X1 U69 ( .A(n103), .ZN(O[31]) );
  AOI22_X1 U70 ( .A1(IN0[31]), .A2(n5), .B1(IN1[31]), .B2(n7), .ZN(n103) );
  INV_X1 U71 ( .A(n99), .ZN(O[28]) );
  AOI22_X1 U72 ( .A1(IN0[28]), .A2(n5), .B1(IN1[28]), .B2(n8), .ZN(n99) );
  INV_X1 U73 ( .A(n100), .ZN(O[29]) );
  AOI22_X1 U74 ( .A1(IN0[29]), .A2(n5), .B1(IN1[29]), .B2(n8), .ZN(n100) );
  INV_X1 U75 ( .A(n79), .ZN(O[0]) );
  AOI22_X1 U76 ( .A1(IN0[0]), .A2(n4), .B1(IN1[0]), .B2(n13), .ZN(n79) );
  INV_X1 U77 ( .A(n101), .ZN(O[2]) );
  INV_X1 U78 ( .A(n105), .ZN(O[4]) );
endmodule


module REG_BITS1 ( CLK, RST, I, O );
  input [0:0] I;
  output [0:0] O;
  input CLK, RST;
  wire   n1;

  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  INV_X1 U2 ( .A(RST), .ZN(n1) );
endmodule


module REG_BITS32_13 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1, n2, n3, n4;

  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n3), .Q(O[31]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n3), .Q(O[30]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n3), .Q(O[29]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n3), .Q(O[28]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n3), .Q(O[26]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n3), .Q(O[25]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n3), .Q(O[24]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n2), .Q(O[23]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n2), .Q(O[22]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n2), .Q(O[21]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n2), .Q(O[20]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n2), .Q(O[19]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n2), .Q(O[18]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n2), .Q(O[17]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n2), .Q(O[16]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n2), .Q(O[15]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n2), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n2), .Q(O[13]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n2), .Q(O[12]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n3), .Q(O[27]) );
  BUF_X1 U2 ( .A(n4), .Z(n1) );
  BUF_X1 U3 ( .A(n4), .Z(n2) );
  BUF_X1 U4 ( .A(n4), .Z(n3) );
  INV_X1 U5 ( .A(RST), .ZN(n4) );
endmodule


module REG_BITS32_12 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1, n2, n3, n4;

  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n3), .Q(O[31]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n3), .Q(O[30]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n3), .Q(O[29]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n3), .Q(O[28]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n3), .Q(O[27]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n3), .Q(O[26]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n3), .Q(O[25]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n3), .Q(O[24]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n2), .Q(O[23]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n2), .Q(O[22]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n2), .Q(O[21]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n2), .Q(O[20]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n2), .Q(O[19]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n2), .Q(O[18]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n2), .Q(O[17]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n2), .Q(O[16]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n2), .Q(O[15]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n2), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n2), .Q(O[13]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n2), .Q(O[12]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  BUF_X1 U2 ( .A(n4), .Z(n1) );
  BUF_X1 U3 ( .A(n4), .Z(n2) );
  BUF_X1 U4 ( .A(n4), .Z(n3) );
  INV_X1 U5 ( .A(RST), .ZN(n4) );
endmodule


module REG_BITS32_11 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1;

  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n1), .Q(O[31]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n1), .Q(O[30]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n1), .Q(O[29]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n1), .Q(O[28]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n1), .Q(O[27]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n1), .Q(O[26]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n1), .Q(O[25]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n1), .Q(O[24]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n1), .Q(O[23]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n1), .Q(O[22]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n1), .Q(O[21]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n1), .Q(O[20]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n1), .Q(O[19]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n1), .Q(O[18]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n1), .Q(O[17]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n1), .Q(O[16]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n1), .Q(O[15]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n1), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n1), .Q(O[13]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n1), .Q(O[12]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  INV_X2 U2 ( .A(RST), .ZN(n1) );
endmodule


module REG_BITS32_10 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1, n2, n3;

  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n2), .Q(O[31]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n2), .Q(O[30]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n2), .Q(O[29]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n2), .Q(O[28]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n3), .Q(O[9]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n3), .Q(O[10]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n3), .Q(O[11]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n3), .Q(O[16]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n3), .Q(O[15]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n3), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n3), .Q(O[13]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n3), .Q(O[17]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n3), .Q(O[12]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n3), .Q(O[6]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n3), .Q(O[8]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n3), .Q(O[26]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n3), .Q(O[5]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n3), .Q(O[2]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n3), .Q(O[27]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n3), .Q(O[25]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n3), .Q(O[4]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n3), .Q(O[21]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n3), .Q(O[3]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n3), .Q(O[7]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n3), .Q(O[23]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n3), .Q(O[22]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n3), .Q(O[24]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n3), .Q(O[20]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n3), .Q(O[18]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n3), .Q(O[19]) );
  INV_X2 U2 ( .A(RST), .ZN(n3) );
  BUF_X1 U3 ( .A(n3), .Z(n1) );
  BUF_X1 U4 ( .A(n3), .Z(n2) );
endmodule


module REG_BITS32_9 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1, n2, n3, n4;

  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n3), .Q(O[31]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n3), .Q(O[30]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n3), .Q(O[29]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n3), .Q(O[28]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n3), .Q(O[27]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n3), .Q(O[26]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n3), .Q(O[25]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n3), .Q(O[24]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n2), .Q(O[23]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n2), .Q(O[22]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n2), .Q(O[21]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n2), .Q(O[20]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n2), .Q(O[19]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n2), .Q(O[18]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n2), .Q(O[17]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n2), .Q(O[16]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n2), .Q(O[15]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n2), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n2), .Q(O[13]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n2), .Q(O[12]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  BUF_X1 U2 ( .A(n4), .Z(n1) );
  BUF_X1 U3 ( .A(n4), .Z(n2) );
  BUF_X1 U4 ( .A(n4), .Z(n3) );
  INV_X1 U5 ( .A(RST), .ZN(n4) );
endmodule


module REG_BITS32_8 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1, n2, n3, n4;

  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n3), .Q(O[31]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n3), .Q(O[30]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n3), .Q(O[29]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n3), .Q(O[28]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n3), .Q(O[27]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n3), .Q(O[26]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n3), .Q(O[25]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n3), .Q(O[24]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n2), .Q(O[23]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n2), .Q(O[22]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n2), .Q(O[21]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n2), .Q(O[20]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n2), .Q(O[19]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n2), .Q(O[18]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n2), .Q(O[17]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n2), .Q(O[16]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n2), .Q(O[15]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n2), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n2), .Q(O[13]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n2), .Q(O[12]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  BUF_X1 U2 ( .A(n4), .Z(n1) );
  BUF_X1 U3 ( .A(n4), .Z(n2) );
  BUF_X1 U4 ( .A(n4), .Z(n3) );
  INV_X1 U5 ( .A(RST), .ZN(n4) );
endmodule


module REG_BITS16 ( CLK, RST, I, O );
  input [15:0] I;
  output [15:0] O;
  input CLK, RST;
  wire   n1;

  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n1), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n1), .Q(O[13]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n1), .Q(O[12]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n1), .Q(O[15]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  INV_X1 U2 ( .A(RST), .ZN(n1) );
endmodule


module REG_BITS5_0 ( CLK, RST, I, O );
  input [4:0] I;
  output [4:0] O;
  input CLK, RST;
  wire   n1;

  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  INV_X1 U2 ( .A(RST), .ZN(n1) );
endmodule


module REG_BITS32_7 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1;

  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n1), .Q(O[31]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n1), .Q(O[27]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n1), .Q(O[23]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n1), .Q(O[30]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n1), .Q(O[29]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n1), .Q(O[28]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n1), .Q(O[26]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n1), .Q(O[25]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n1), .Q(O[24]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n1), .Q(O[22]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n1), .Q(O[21]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n1), .Q(O[20]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n1), .Q(O[19]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n1), .Q(O[18]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n1), .Q(O[17]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n1), .Q(O[16]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n1), .Q(O[15]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n1), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n1), .Q(O[13]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n1), .Q(O[12]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  INV_X2 U2 ( .A(RST), .ZN(n1) );
endmodule


module REG_BITS32_6 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1;

  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n1), .Q(O[16]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n1), .Q(O[12]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n1), .Q(O[17]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n1), .Q(O[20]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n1), .Q(O[13]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n1), .Q(O[18]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n1), .Q(O[24]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n1), .Q(O[21]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n1), .Q(O[19]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n1), .Q(O[14]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n1), .Q(O[22]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n1), .Q(O[25]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n1), .Q(O[15]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n1), .Q(O[28]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n1), .Q(O[23]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n1), .Q(O[26]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n1), .Q(O[27]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n1), .Q(O[29]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n1), .Q(O[30]) );
  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n1), .Q(O[31]) );
  INV_X2 U2 ( .A(RST), .ZN(n1) );
endmodule


module REG_BITS32_5 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1;

  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n1), .Q(O[16]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n1), .Q(O[18]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n1), .Q(O[20]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n1), .Q(O[17]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n1), .Q(O[12]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n1), .Q(O[21]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n1), .Q(O[19]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n1), .Q(O[22]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n1), .Q(O[24]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n1), .Q(O[13]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n1), .Q(O[14]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n1), .Q(O[25]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n1), .Q(O[26]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n1), .Q(O[28]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n1), .Q(O[23]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n1), .Q(O[29]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n1), .Q(O[15]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n1), .Q(O[30]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n1), .Q(O[27]) );
  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n1), .Q(O[31]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  INV_X2 U2 ( .A(RST), .ZN(n1) );
endmodule


module REG_BITS32_4 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1;

  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n1), .Q(O[19]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n1), .Q(O[18]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n1), .Q(O[17]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n1), .Q(O[16]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n1), .Q(O[15]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n1), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n1), .Q(O[13]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n1), .Q(O[12]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n1), .Q(O[31]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n1), .Q(O[30]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n1), .Q(O[29]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n1), .Q(O[28]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n1), .Q(O[27]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n1), .Q(O[26]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n1), .Q(O[25]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n1), .Q(O[24]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n1), .Q(O[23]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n1), .Q(O[22]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n1), .Q(O[21]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n1), .Q(O[20]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  INV_X2 U2 ( .A(RST), .ZN(n1) );
endmodule


module REG_BITS5_2 ( CLK, RST, I, O );
  input [4:0] I;
  output [4:0] O;
  input CLK, RST;
  wire   n1;

  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  INV_X1 U2 ( .A(RST), .ZN(n1) );
endmodule


module REG_BITS32_3 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1;

  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n1), .Q(O[31]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n1), .Q(O[30]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n1), .Q(O[29]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n1), .Q(O[28]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n1), .Q(O[27]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n1), .Q(O[26]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n1), .Q(O[25]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n1), .Q(O[24]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n1), .Q(O[23]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n1), .Q(O[22]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n1), .Q(O[21]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n1), .Q(O[20]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n1), .Q(O[19]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n1), .Q(O[18]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n1), .Q(O[17]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n1), .Q(O[16]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n1), .Q(O[15]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n1), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n1), .Q(O[13]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n1), .Q(O[12]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  INV_X2 U2 ( .A(RST), .ZN(n1) );
endmodule


module REG_BITS32_2 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1, n2, n3, n4;

  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n3), .Q(O[31]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n3), .Q(O[30]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n3), .Q(O[29]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n3), .Q(O[28]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n3), .Q(O[27]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n3), .Q(O[26]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n3), .Q(O[25]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n3), .Q(O[24]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n2), .Q(O[23]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n2), .Q(O[22]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n2), .Q(O[21]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n2), .Q(O[20]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n2), .Q(O[19]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n2), .Q(O[18]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n2), .Q(O[17]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n2), .Q(O[16]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n2), .Q(O[15]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n2), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n2), .Q(O[13]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n2), .Q(O[12]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  BUF_X1 U2 ( .A(n4), .Z(n1) );
  BUF_X1 U3 ( .A(n4), .Z(n2) );
  BUF_X1 U4 ( .A(n4), .Z(n3) );
  INV_X1 U5 ( .A(RST), .ZN(n4) );
endmodule


module REG_BITS32_1 ( CLK, RST, I, O );
  input [31:0] I;
  output [31:0] O;
  input CLK, RST;
  wire   n1;

  DFFR_X1 \O_reg[31]  ( .D(I[31]), .CK(CLK), .RN(n1), .Q(O[31]) );
  DFFR_X1 \O_reg[30]  ( .D(I[30]), .CK(CLK), .RN(n1), .Q(O[30]) );
  DFFR_X1 \O_reg[29]  ( .D(I[29]), .CK(CLK), .RN(n1), .Q(O[29]) );
  DFFR_X1 \O_reg[28]  ( .D(I[28]), .CK(CLK), .RN(n1), .Q(O[28]) );
  DFFR_X1 \O_reg[27]  ( .D(I[27]), .CK(CLK), .RN(n1), .Q(O[27]) );
  DFFR_X1 \O_reg[26]  ( .D(I[26]), .CK(CLK), .RN(n1), .Q(O[26]) );
  DFFR_X1 \O_reg[25]  ( .D(I[25]), .CK(CLK), .RN(n1), .Q(O[25]) );
  DFFR_X1 \O_reg[24]  ( .D(I[24]), .CK(CLK), .RN(n1), .Q(O[24]) );
  DFFR_X1 \O_reg[23]  ( .D(I[23]), .CK(CLK), .RN(n1), .Q(O[23]) );
  DFFR_X1 \O_reg[22]  ( .D(I[22]), .CK(CLK), .RN(n1), .Q(O[22]) );
  DFFR_X1 \O_reg[21]  ( .D(I[21]), .CK(CLK), .RN(n1), .Q(O[21]) );
  DFFR_X1 \O_reg[20]  ( .D(I[20]), .CK(CLK), .RN(n1), .Q(O[20]) );
  DFFR_X1 \O_reg[19]  ( .D(I[19]), .CK(CLK), .RN(n1), .Q(O[19]) );
  DFFR_X1 \O_reg[18]  ( .D(I[18]), .CK(CLK), .RN(n1), .Q(O[18]) );
  DFFR_X1 \O_reg[17]  ( .D(I[17]), .CK(CLK), .RN(n1), .Q(O[17]) );
  DFFR_X1 \O_reg[16]  ( .D(I[16]), .CK(CLK), .RN(n1), .Q(O[16]) );
  DFFR_X1 \O_reg[15]  ( .D(I[15]), .CK(CLK), .RN(n1), .Q(O[15]) );
  DFFR_X1 \O_reg[14]  ( .D(I[14]), .CK(CLK), .RN(n1), .Q(O[14]) );
  DFFR_X1 \O_reg[13]  ( .D(I[13]), .CK(CLK), .RN(n1), .Q(O[13]) );
  DFFR_X1 \O_reg[12]  ( .D(I[12]), .CK(CLK), .RN(n1), .Q(O[12]) );
  DFFR_X1 \O_reg[11]  ( .D(I[11]), .CK(CLK), .RN(n1), .Q(O[11]) );
  DFFR_X1 \O_reg[10]  ( .D(I[10]), .CK(CLK), .RN(n1), .Q(O[10]) );
  DFFR_X1 \O_reg[9]  ( .D(I[9]), .CK(CLK), .RN(n1), .Q(O[9]) );
  DFFR_X1 \O_reg[8]  ( .D(I[8]), .CK(CLK), .RN(n1), .Q(O[8]) );
  DFFR_X1 \O_reg[7]  ( .D(I[7]), .CK(CLK), .RN(n1), .Q(O[7]) );
  DFFR_X1 \O_reg[6]  ( .D(I[6]), .CK(CLK), .RN(n1), .Q(O[6]) );
  DFFR_X1 \O_reg[5]  ( .D(I[5]), .CK(CLK), .RN(n1), .Q(O[5]) );
  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  INV_X2 U2 ( .A(RST), .ZN(n1) );
endmodule


module REG_BITS5_1 ( CLK, RST, I, O );
  input [4:0] I;
  output [4:0] O;
  input CLK, RST;
  wire   n1;

  DFFR_X1 \O_reg[4]  ( .D(I[4]), .CK(CLK), .RN(n1), .Q(O[4]) );
  DFFR_X1 \O_reg[3]  ( .D(I[3]), .CK(CLK), .RN(n1), .Q(O[3]) );
  DFFR_X1 \O_reg[2]  ( .D(I[2]), .CK(CLK), .RN(n1), .Q(O[2]) );
  DFFR_X1 \O_reg[1]  ( .D(I[1]), .CK(CLK), .RN(n1), .Q(O[1]) );
  DFFR_X1 \O_reg[0]  ( .D(I[0]), .CK(CLK), .RN(n1), .Q(O[0]) );
  INV_X1 U2 ( .A(RST), .ZN(n1) );
endmodule


module DP ( CLK, RST, INSTRUCTION, DATA_IN, RegDst, RegWrite, ALUSrc, 
        ALUOpcode, MemToReg, Jump, Branch, Jal, PC_OUT, ALU_OUT, DATA_OUT, 
        INSTRUCTION_IF_ID_OUT );
  input [31:0] INSTRUCTION;
  input [31:0] DATA_IN;
  input [3:0] ALUOpcode;
  output [31:0] PC_OUT;
  output [31:0] ALU_OUT;
  output [31:0] DATA_OUT;
  output [31:0] INSTRUCTION_IF_ID_OUT;
  input CLK, RST, RegDst, RegWrite, ALUSrc, MemToReg, Jump, Branch, Jal;
  wire   ZERO_i, SE_SEL_i, \PC_MUX_SEL_i[0] , n3, n1, n2, n4, n5, n6, n7, n8,
         n9, n10, n11;
  wire   [15:0] SE_IMM_i;
  wire   [31:0] PC_IN_i;
  wire   [31:0] PC_ADDER_OUT_i;
  wire   [4:0] ADDR_WR_MUX_OUT_i;
  wire   [31:0] MEM_MUX_OUT_i;
  wire   [31:0] PC_ADDER_REG_MEM_WB_i;
  wire   [31:0] JAL_MUX_OUT_i;
  wire   [4:0] ADDR_WR_MUX_OUT_REG_MEM_WB_i;
  wire   [4:0] JAL_R31_ADDR_MUX_OUT_i;
  wire   [31:0] DATA_OUT1_i;
  wire   [31:0] DATA_OUT2_i;
  wire   [31:0] RF_DATA_OUT2_REG_ID_EX_i;
  wire   [31:0] SE_OUT_MUX_i;
  wire   [31:0] ALU_MUX_OUT_i;
  wire   [31:0] RF_DATA_OUT1_REG_ID_EX_i;
  wire   [31:0] ALU_OUT_i;
  wire   [31:0] JLABEL_REG_ID_EX_i;
  wire   [31:0] PC_OFFSET_i;
  wire   [31:0] PC_ADDER_REG_ID_EX_i;
  wire   [31:0] PC_BRANCH_ADDER_OUT_i;
  wire   [31:0] PC_BRANCH_ADDER_OUT_REG_EX_MEM_i;
  wire   [31:0] ALU_OUT_REG_MEM_WB_i;
  wire   [31:0] DATA_IN_REG_MEM_WB_i;
  wire   [31:0] PC_ADDER_REG_IF_ID_i;
  wire   [4:0] ADDR_WR_MUX_OUT_REG_ID_EX_i;
  wire   [31:0] PC_ADDER_REG_EX_MEM_i;
  wire   [4:0] ADDR_WR_MUX_OUT_REG_EX_MEM_i;

  REG_BITS32_0 PC ( .CLK(n11), .RST(n9), .I(PC_IN_i), .O(PC_OUT) );
  ADDER_0 PC_ADDER ( .A(PC_OUT), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b0}), .S(PC_ADDER_OUT_i) );
  MUX21_NBIT5_0 ADDR_WR_MUX ( .IN0(INSTRUCTION_IF_ID_OUT[20:16]), .IN1(
        INSTRUCTION_IF_ID_OUT[15:11]), .S(RegDst), .O(ADDR_WR_MUX_OUT_i) );
  MUX21_NBIT32_0 JAL_MUX ( .IN0(MEM_MUX_OUT_i), .IN1(PC_ADDER_REG_MEM_WB_i), 
        .S(Jal), .O(JAL_MUX_OUT_i) );
  MUX21_NBIT5_1 JAL_R31_ADDR ( .IN0(ADDR_WR_MUX_OUT_REG_MEM_WB_i), .IN1({1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .S(Jal), .O(JAL_R31_ADDR_MUX_OUT_i) );
  RF REGFILE ( .RST(n7), .WE(RegWrite), .ADDR_RD1(INSTRUCTION_IF_ID_OUT[25:21]), .ADDR_RD2(INSTRUCTION_IF_ID_OUT[20:16]), .ADDR_WR(JAL_R31_ADDR_MUX_OUT_i), 
        .DATA_IN(JAL_MUX_OUT_i), .DATA_OUT1(DATA_OUT1_i), .DATA_OUT2(
        DATA_OUT2_i) );
  MUX21_NBIT32_5 ALU_MUX ( .IN0(RF_DATA_OUT2_REG_ID_EX_i), .IN1(SE_OUT_MUX_i), 
        .S(ALUSrc), .O(ALU_MUX_OUT_i) );
  ALU ALU_DP ( .OP1(RF_DATA_OUT1_REG_ID_EX_i), .OP2(ALU_MUX_OUT_i), .ALU_OP(
        ALUOpcode), .RES(ALU_OUT_i), .ZERO(ZERO_i) );
  MUX21_NBIT32_4 JUMP_MUX ( .IN0(JLABEL_REG_ID_EX_i), .IN1({n5, n5, n5, n5, n5, 
        n5, n6, n6, n6, n6, n6, n6, n6, n6, n6, n6, n6, SE_IMM_i[14:0]}), .S(
        n10), .O(PC_OFFSET_i) );
  ADDER_1 PC_BRANCH_ADDER ( .A(PC_ADDER_REG_ID_EX_i), .B(PC_OFFSET_i), .S(
        PC_BRANCH_ADDER_OUT_i) );
  MUX21_NBIT32_3 PC_MUX ( .IN0({n2, PC_ADDER_OUT_i[30:28], n1, 
        PC_ADDER_OUT_i[26:0]}), .IN1(PC_BRANCH_ADDER_OUT_REG_EX_MEM_i), .S(
        \PC_MUX_SEL_i[0] ), .O(PC_IN_i) );
  MUX21_NBIT32_2 MEM_MUX ( .IN0(ALU_OUT_REG_MEM_WB_i), .IN1(
        DATA_IN_REG_MEM_WB_i), .S(MemToReg), .O(MEM_MUX_OUT_i) );
  MUX21_NBIT32_1 SE_MUX ( .IN0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n4, SE_IMM_i[14:0]}), 
        .IN1({n4, n4, n4, n4, n4, n4, n4, n4, n4, n4, n4, n5, n5, n5, n5, n5, 
        n5, SE_IMM_i[14:0]}), .S(SE_SEL_i), .O(SE_OUT_MUX_i) );
  REG_BITS1 PC_SRC_EX_MEM ( .CLK(CLK), .RST(n9), .I(n10), .O(\PC_MUX_SEL_i[0] ) );
  REG_BITS32_13 PC_ADDER_REG_IF_ID ( .CLK(CLK), .RST(n9), .I(PC_ADDER_OUT_i), 
        .O(PC_ADDER_REG_IF_ID_i) );
  REG_BITS32_12 INSTRMEM_REG_IF_ID ( .CLK(CLK), .RST(n9), .I(INSTRUCTION), .O(
        INSTRUCTION_IF_ID_OUT) );
  REG_BITS32_11 PC_ADDER_REG_ID_EX ( .CLK(CLK), .RST(n8), .I(
        PC_ADDER_REG_IF_ID_i), .O(PC_ADDER_REG_ID_EX_i) );
  REG_BITS32_10 JLABEL_REG_ID_EX ( .CLK(CLK), .RST(n9), .I({1'b0, 1'b0, 1'b0, 
        1'b0, INSTRUCTION_IF_ID_OUT[25:0], 1'b0, 1'b0}), .O(JLABEL_REG_ID_EX_i) );
  REG_BITS32_9 RF_DATA_OUT1_REG_ID_EX ( .CLK(CLK), .RST(n8), .I(DATA_OUT1_i), 
        .O(RF_DATA_OUT1_REG_ID_EX_i) );
  REG_BITS32_8 RF_DATA_OUT2_REG_ID_EX ( .CLK(CLK), .RST(n8), .I(DATA_OUT2_i), 
        .O(RF_DATA_OUT2_REG_ID_EX_i) );
  REG_BITS16 IMM_REG_ID_EX ( .CLK(CLK), .RST(n9), .I(
        INSTRUCTION_IF_ID_OUT[15:0]), .O(SE_IMM_i) );
  REG_BITS5_0 ADDR_WR_MUX_OUT_REG_ID_EX ( .CLK(CLK), .RST(n7), .I(
        ADDR_WR_MUX_OUT_i), .O(ADDR_WR_MUX_OUT_REG_ID_EX_i) );
  REG_BITS32_7 PC_ADDER_REG_EX_MEM ( .CLK(CLK), .RST(n8), .I(
        PC_ADDER_REG_ID_EX_i), .O(PC_ADDER_REG_EX_MEM_i) );
  REG_BITS32_6 PC_BRANCH_ADDER_OUT_REG_EX_MEM ( .CLK(CLK), .RST(n8), .I(
        PC_BRANCH_ADDER_OUT_i), .O(PC_BRANCH_ADDER_OUT_REG_EX_MEM_i) );
  REG_BITS32_5 ALU_OUT_REG_EX_MEM ( .CLK(CLK), .RST(n8), .I(ALU_OUT_i), .O(
        ALU_OUT) );
  REG_BITS32_4 RF_DATA_OUT2_REG_EX_MEM ( .CLK(CLK), .RST(n7), .I(
        RF_DATA_OUT2_REG_ID_EX_i), .O(DATA_OUT) );
  REG_BITS5_2 ADDR_WR_MUX_OUT_REG_EX_MEM ( .CLK(CLK), .RST(n9), .I(
        ADDR_WR_MUX_OUT_REG_ID_EX_i), .O(ADDR_WR_MUX_OUT_REG_EX_MEM_i) );
  REG_BITS32_3 PC_ADDER_REG_MEM_WB ( .CLK(CLK), .RST(n7), .I(
        PC_ADDER_REG_EX_MEM_i), .O(PC_ADDER_REG_MEM_WB_i) );
  REG_BITS32_2 DATA_IN_REG_MEM_WB ( .CLK(CLK), .RST(n7), .I(DATA_IN), .O(
        DATA_IN_REG_MEM_WB_i) );
  REG_BITS32_1 ALU_OUT_REG_MEM_WB ( .CLK(CLK), .RST(n7), .I(ALU_OUT), .O(
        ALU_OUT_REG_MEM_WB_i) );
  REG_BITS5_1 ADDR_WR_MUX_OUT_REG_MEM_WB ( .CLK(CLK), .RST(n9), .I(
        ADDR_WR_MUX_OUT_REG_EX_MEM_i), .O(ADDR_WR_MUX_OUT_REG_MEM_WB_i) );
  BUF_X1 U3 ( .A(RST), .Z(n9) );
  CLKBUF_X1 U4 ( .A(PC_ADDER_OUT_i[27]), .Z(n1) );
  BUF_X1 U5 ( .A(SE_IMM_i[15]), .Z(n4) );
  BUF_X1 U6 ( .A(SE_IMM_i[15]), .Z(n5) );
  BUF_X1 U7 ( .A(SE_IMM_i[15]), .Z(n6) );
  NOR2_X1 U8 ( .A1(ALUOpcode[3]), .A2(ALUOpcode[2]), .ZN(SE_SEL_i) );
  INV_X1 U9 ( .A(n3), .ZN(n10) );
  AOI21_X1 U10 ( .B1(ZERO_i), .B2(Branch), .A(Jump), .ZN(n3) );
  INV_X1 U11 ( .A(CLK), .ZN(n11) );
  CLKBUF_X1 U12 ( .A(PC_ADDER_OUT_i[31]), .Z(n2) );
  CLKBUF_X1 U13 ( .A(RST), .Z(n7) );
  CLKBUF_X1 U14 ( .A(RST), .Z(n8) );
endmodule


module HWCU ( OPCODE, FUNC, CLK, RST, ALUSrc, Jump, Branch, ALUOpcode, WE, RE, 
        MemToReg, RegDst, Jal, RegWrite );
  input [5:0] OPCODE;
  input [10:0] FUNC;
  output [3:0] ALUOpcode;
  input CLK, RST;
  output ALUSrc, Jump, Branch, WE, RE, MemToReg, RegDst, Jal, RegWrite;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20;
  wire   [3:0] next_aluopcode;
  assign ALUSrc = 1'b0;
  assign Jump = 1'b0;
  assign Branch = 1'b0;
  assign WE = 1'b0;
  assign RE = 1'b0;
  assign MemToReg = 1'b0;
  assign Jal = 1'b0;
  assign RegWrite = 1'b0;
  assign RegDst = 1'b0;

  OAI33_X1 U58 ( .A1(n23), .A2(FUNC[2]), .A3(n24), .B1(n25), .B2(n26), .B3(n27), .ZN(n22) );
  NAND3_X1 U59 ( .A1(n16), .A2(n15), .A3(n28), .ZN(n25) );
  NAND3_X1 U60 ( .A1(n32), .A2(n9), .A3(OPCODE[3]), .ZN(n30) );
  NAND3_X1 U61 ( .A1(n3), .A2(n29), .A3(n37), .ZN(next_aluopcode[1]) );
  OAI33_X1 U62 ( .A1(n36), .A2(OPCODE[0]), .A3(n10), .B1(n40), .B2(n8), .B3(n7), .ZN(n39) );
  NAND3_X1 U63 ( .A1(n4), .A2(n3), .A3(n44), .ZN(next_aluopcode[0]) );
  NAND3_X1 U64 ( .A1(n42), .A2(n9), .A3(OPCODE[1]), .ZN(n48) );
  NAND3_X1 U65 ( .A1(n50), .A2(n17), .A3(n19), .ZN(n49) );
  NAND3_X1 U66 ( .A1(n28), .A2(n16), .A3(FUNC[5]), .ZN(n33) );
  OAI33_X1 U67 ( .A1(n7), .A2(OPCODE[0]), .A3(n6), .B1(n52), .B2(n13), .B3(n27), .ZN(n51) );
  NAND3_X1 U68 ( .A1(FUNC[3]), .A2(n28), .A3(FUNC[5]), .ZN(n24) );
  NAND3_X1 U69 ( .A1(n50), .A2(n18), .A3(FUNC[0]), .ZN(n23) );
  DFFR_X1 \curr_aluopcode_reg[3]  ( .D(next_aluopcode[3]), .CK(CLK), .RN(n1), 
        .Q(ALUOpcode[3]) );
  DFFR_X1 \curr_aluopcode_reg[0]  ( .D(next_aluopcode[0]), .CK(CLK), .RN(n1), 
        .Q(ALUOpcode[0]) );
  DFFR_X1 \curr_aluopcode_reg[2]  ( .D(next_aluopcode[2]), .CK(CLK), .RN(n1), 
        .Q(ALUOpcode[2]) );
  DFFR_X1 \curr_aluopcode_reg[1]  ( .D(next_aluopcode[1]), .CK(CLK), .RN(n1), 
        .Q(ALUOpcode[1]) );
  OAI221_X1 U11 ( .B1(n33), .B2(n34), .C1(n35), .C2(n36), .A(n3), .ZN(
        next_aluopcode[2]) );
  NOR2_X1 U12 ( .A1(n12), .A2(n10), .ZN(n35) );
  OAI21_X1 U13 ( .B1(n18), .B2(n20), .A(n2), .ZN(n34) );
  AOI21_X1 U14 ( .B1(n41), .B2(n42), .A(n43), .ZN(n29) );
  INV_X1 U15 ( .A(n41), .ZN(n6) );
  INV_X1 U16 ( .A(n33), .ZN(n14) );
  INV_X1 U17 ( .A(n27), .ZN(n2) );
  INV_X1 U18 ( .A(n53), .ZN(n4) );
  AOI211_X1 U19 ( .C1(n14), .C2(n45), .A(n43), .B(n46), .ZN(n44) );
  OAI22_X1 U20 ( .A1(n23), .A2(n24), .B1(n36), .B2(n11), .ZN(n53) );
  INV_X1 U21 ( .A(n32), .ZN(n11) );
  NOR4_X1 U22 ( .A1(FUNC[6]), .A2(FUNC[4]), .A3(FUNC[10]), .A4(n54), .ZN(n28)
         );
  OR3_X1 U23 ( .A1(FUNC[9]), .A2(FUNC[8]), .A3(FUNC[7]), .ZN(n54) );
  NOR4_X1 U24 ( .A1(n9), .A2(OPCODE[1]), .A3(OPCODE[3]), .A4(OPCODE[5]), .ZN(
        n41) );
  NOR3_X1 U25 ( .A1(n6), .A2(OPCODE[4]), .A3(n12), .ZN(n43) );
  AOI211_X1 U26 ( .C1(n47), .C2(n48), .A(n8), .B(OPCODE[5]), .ZN(n46) );
  NAND2_X1 U27 ( .A1(OPCODE[4]), .A2(n32), .ZN(n47) );
  NOR2_X1 U28 ( .A1(n12), .A2(OPCODE[1]), .ZN(n32) );
  NOR2_X1 U29 ( .A1(OPCODE[0]), .A2(OPCODE[4]), .ZN(n42) );
  NAND4_X1 U30 ( .A1(OPCODE[1]), .A2(OPCODE[2]), .A3(n12), .A4(n8), .ZN(n31)
         );
  INV_X1 U31 ( .A(OPCODE[2]), .ZN(n9) );
  OAI21_X1 U32 ( .B1(n17), .B2(n23), .A(n49), .ZN(n45) );
  INV_X1 U33 ( .A(FUNC[2]), .ZN(n17) );
  INV_X1 U34 ( .A(n26), .ZN(n19) );
  OR4_X1 U35 ( .A1(n8), .A2(n9), .A3(OPCODE[4]), .A4(OPCODE[5]), .ZN(n36) );
  INV_X1 U36 ( .A(OPCODE[0]), .ZN(n12) );
  INV_X1 U37 ( .A(n51), .ZN(n3) );
  NAND4_X1 U38 ( .A1(n20), .A2(n18), .A3(n16), .A4(n15), .ZN(n52) );
  INV_X1 U39 ( .A(n28), .ZN(n13) );
  INV_X1 U40 ( .A(OPCODE[3]), .ZN(n8) );
  NAND2_X1 U41 ( .A1(FUNC[1]), .A2(n20), .ZN(n26) );
  INV_X1 U42 ( .A(OPCODE[1]), .ZN(n10) );
  INV_X1 U43 ( .A(FUNC[0]), .ZN(n20) );
  NAND2_X1 U44 ( .A1(FUNC[2]), .A2(n50), .ZN(n27) );
  INV_X1 U45 ( .A(FUNC[1]), .ZN(n18) );
  INV_X1 U46 ( .A(OPCODE[4]), .ZN(n7) );
  AND4_X1 U47 ( .A1(n42), .A2(n10), .A3(n55), .A4(n9), .ZN(n50) );
  NOR2_X1 U48 ( .A1(OPCODE[5]), .A2(OPCODE[3]), .ZN(n55) );
  INV_X1 U49 ( .A(FUNC[3]), .ZN(n16) );
  AOI21_X1 U50 ( .B1(n2), .B2(n38), .A(n39), .ZN(n37) );
  OAI22_X1 U51 ( .A1(FUNC[1]), .A2(n24), .B1(n26), .B2(n33), .ZN(n38) );
  INV_X1 U52 ( .A(FUNC[5]), .ZN(n15) );
  OR3_X1 U53 ( .A1(OPCODE[1]), .A2(OPCODE[5]), .A3(n9), .ZN(n40) );
  OR3_X1 U54 ( .A1(n21), .A2(n5), .A3(n22), .ZN(next_aluopcode[3]) );
  AOI211_X1 U55 ( .C1(n30), .C2(n31), .A(n7), .B(OPCODE[5]), .ZN(n21) );
  INV_X1 U56 ( .A(n29), .ZN(n5) );
  INV_X1 U57 ( .A(RST), .ZN(n1) );
endmodule


module CPU ( CLK, RST );
  input CLK, RST;
  wire   INSTR_IF_ID_i_31, INSTR_IF_ID_i_30, INSTR_IF_ID_i_29,
         INSTR_IF_ID_i_28, INSTR_IF_ID_i_27, INSTR_IF_ID_i_26;
  wire   [31:0] INSTR_i;
  wire   [31:0] DATA_IN_i;
  wire   [3:0] ALUOpcode_i;
  wire   [31:0] PC_OUT_i;
  wire   [31:0] ALU_OUT_i;
  wire   [31:0] DATA_OUT_i;
  wire   [10:0] INSTR_IF_ID_i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14;

  DP CPU_DP ( .CLK(CLK), .RST(RST), .INSTRUCTION(INSTR_i), .DATA_IN(DATA_IN_i), 
        .RegDst(1'b0), .RegWrite(1'b0), .ALUSrc(1'b0), .ALUOpcode(ALUOpcode_i), 
        .MemToReg(1'b0), .Jump(1'b0), .Branch(1'b0), .Jal(1'b0), .PC_OUT(
        PC_OUT_i), .ALU_OUT(ALU_OUT_i), .DATA_OUT(DATA_OUT_i), 
        .INSTRUCTION_IF_ID_OUT({INSTR_IF_ID_i_31, INSTR_IF_ID_i_30, 
        INSTR_IF_ID_i_29, INSTR_IF_ID_i_28, INSTR_IF_ID_i_27, INSTR_IF_ID_i_26, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, INSTR_IF_ID_i}) );
  INSTRMEM CPU_INSTRMEM ( .ADDR_RD(PC_OUT_i), .DATA_OUT(INSTR_i) );
  DATAMEM CPU_DATAMEM ( .RST(RST), .RE(1'b0), .WE(1'b0), .ADDR(ALU_OUT_i), 
        .DATA_IN(DATA_OUT_i), .DATA_OUT(DATA_IN_i) );
  HWCU CPU_CU ( .OPCODE({INSTR_IF_ID_i_31, INSTR_IF_ID_i_30, INSTR_IF_ID_i_29, 
        INSTR_IF_ID_i_28, INSTR_IF_ID_i_27, INSTR_IF_ID_i_26}), .FUNC(
        INSTR_IF_ID_i), .CLK(CLK), .RST(RST), .ALUOpcode(ALUOpcode_i) );
endmodule

